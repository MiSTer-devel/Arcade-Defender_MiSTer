library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity defender_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of defender_prog is
	type rom is array(0 to  26623) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"4A",X"DE",X"63",X"A7",X"44",X"AF",X"42",X"7E",X"E8",X"56",X"9E",X"63",X"8D",X"07",X"33",X"84",
		X"7E",X"E8",X"56",X"AE",X"06",X"34",X"46",X"CE",X"A0",X"5F",X"AC",X"C4",X"26",X"18",X"EC",X"84",
		X"ED",X"C4",X"A6",X"06",X"27",X"06",X"DC",X"69",X"9F",X"69",X"20",X"04",X"DC",X"61",X"9F",X"61",
		X"ED",X"84",X"30",X"C4",X"35",X"C6",X"EE",X"C4",X"26",X"E0",X"12",X"7E",X"D7",X"38",X"34",X"62",
		X"DE",X"69",X"26",X"01",X"BD",X"D0",X"3A",X"10",X"AE",X"C4",X"10",X"9F",X"69",X"86",X"01",X"A7",
		X"46",X"A6",X"E4",X"20",X"11",X"34",X"62",X"DE",X"61",X"26",X"03",X"BD",X"D0",X"3A",X"10",X"AE",
		X"C4",X"10",X"9F",X"61",X"6F",X"46",X"AF",X"42",X"A7",X"45",X"86",X"01",X"A7",X"44",X"AE",X"9F",
		X"A0",X"63",X"EF",X"9F",X"A0",X"63",X"AF",X"C4",X"30",X"C4",X"35",X"E2",X"34",X"12",X"8E",X"A0",
		X"5F",X"AE",X"84",X"27",X"0E",X"9C",X"63",X"27",X"F8",X"A6",X"05",X"81",X"02",X"27",X"F2",X"8D",
		X"84",X"20",X"EE",X"35",X"92",X"8D",X"16",X"34",X"66",X"EF",X"06",X"EE",X"66",X"37",X"26",X"ED",
		X"02",X"10",X"AF",X"08",X"37",X"06",X"ED",X"88",X"12",X"EF",X"66",X"35",X"E6",X"34",X"46",X"9E",
		X"67",X"26",X"03",X"BD",X"D0",X"3A",X"EC",X"84",X"DD",X"67",X"DC",X"65",X"ED",X"84",X"4F",X"5F",
		X"ED",X"04",X"A7",X"88",X"14",X"35",X"C6",X"34",X"70",X"CE",X"A0",X"65",X"AC",X"C4",X"26",X"10",
		X"10",X"AE",X"D4",X"10",X"AF",X"C4",X"10",X"9E",X"67",X"9F",X"67",X"10",X"AF",X"84",X"35",X"F0",
		X"EE",X"C4",X"26",X"E8",X"CE",X"A0",X"6B",X"AC",X"C4",X"27",X"E5",X"EE",X"C4",X"26",X"F8",X"BD",
		X"D0",X"3A",X"34",X"70",X"CE",X"A0",X"6D",X"20",X"EE",X"34",X"18",X"10",X"DF",X"77",X"24",X"02",
		X"31",X"22",X"10",X"EE",X"22",X"CB",X"08",X"1F",X"03",X"20",X"4E",X"34",X"18",X"CB",X"08",X"1F",
		X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"1F",X"8B",X"1C",X"00",X"20",X"6A",X"34",
		X"18",X"CB",X"08",X"1F",X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"1F",X"8B",X"1C",
		X"00",X"36",X"3F",X"33",X"C9",X"01",X"08",X"20",X"44",X"34",X"18",X"10",X"DF",X"77",X"24",X"02",
		X"31",X"22",X"10",X"EE",X"22",X"CB",X"08",X"1F",X"03",X"35",X"3F",X"36",X"3F",X"33",X"C9",X"01",
		X"08",X"35",X"3F",X"36",X"3F",X"33",X"C9",X"01",X"08",X"35",X"3F",X"36",X"3F",X"33",X"C9",X"01",
		X"08",X"35",X"3F",X"36",X"3F",X"10",X"FE",X"A0",X"77",X"35",X"98",X"34",X"18",X"CB",X"08",X"1F",
		X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"1F",X"8B",X"1C",X"00",X"36",X"3F",X"33",
		X"C9",X"01",X"08",X"36",X"3F",X"33",X"C9",X"01",X"08",X"36",X"3F",X"33",X"C9",X"01",X"08",X"36",
		X"3F",X"35",X"98",X"34",X"18",X"10",X"DF",X"77",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",
		X"08",X"1F",X"03",X"35",X"3F",X"36",X"3F",X"33",X"C9",X"01",X"08",X"20",X"9C",X"24",X"02",X"31",
		X"22",X"10",X"AE",X"22",X"1F",X"03",X"EC",X"A4",X"ED",X"C4",X"EC",X"22",X"ED",X"42",X"EC",X"24",
		X"ED",X"C9",X"01",X"00",X"EC",X"26",X"ED",X"C9",X"01",X"02",X"EC",X"28",X"ED",X"C9",X"02",X"00",
		X"EC",X"2A",X"ED",X"C9",X"02",X"02",X"39",X"1F",X"03",X"CC",X"00",X"00",X"ED",X"C4",X"ED",X"42",
		X"ED",X"C9",X"01",X"00",X"ED",X"C9",X"01",X"02",X"ED",X"C9",X"02",X"00",X"ED",X"C9",X"02",X"02",
		X"39",X"24",X"02",X"31",X"22",X"10",X"AE",X"22",X"1F",X"03",X"EC",X"A4",X"ED",X"C4",X"EC",X"22",
		X"A7",X"42",X"E7",X"C9",X"01",X"00",X"EC",X"24",X"ED",X"C9",X"01",X"01",X"39",X"1F",X"03",X"CC",
		X"00",X"00",X"ED",X"C4",X"A7",X"42",X"ED",X"C9",X"01",X"00",X"A7",X"C9",X"01",X"02",X"39",X"34",
		X"56",X"10",X"DF",X"77",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"04",X"1F",X"03",X"35",
		X"16",X"36",X"16",X"33",X"C9",X"01",X"04",X"35",X"16",X"36",X"16",X"33",X"C9",X"01",X"04",X"35",
		X"16",X"36",X"16",X"33",X"C9",X"01",X"04",X"35",X"16",X"36",X"16",X"33",X"C9",X"01",X"04",X"35",
		X"16",X"36",X"16",X"33",X"C9",X"01",X"04",X"35",X"16",X"36",X"16",X"10",X"DE",X"77",X"35",X"D6",
		X"34",X"56",X"CB",X"04",X"1F",X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"36",X"16",X"33",X"C9",
		X"01",X"04",X"36",X"16",X"33",X"C9",X"01",X"04",X"36",X"16",X"33",X"C9",X"01",X"04",X"36",X"16",
		X"33",X"C9",X"01",X"04",X"36",X"16",X"33",X"C9",X"01",X"04",X"36",X"16",X"35",X"D6",X"34",X"10",
		X"10",X"DF",X"77",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"06",X"1F",X"03",X"35",X"36",
		X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",
		X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",
		X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",
		X"36",X"36",X"33",X"C9",X"01",X"06",X"35",X"36",X"36",X"36",X"10",X"DE",X"77",X"35",X"90",X"34",
		X"10",X"CB",X"06",X"1F",X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"36",X"36",X"33",
		X"C9",X"01",X"06",X"36",X"36",X"33",X"C9",X"01",X"06",X"36",X"36",X"33",X"C9",X"01",X"06",X"36",
		X"36",X"33",X"C9",X"01",X"06",X"36",X"36",X"33",X"C9",X"01",X"06",X"36",X"36",X"33",X"C9",X"01",
		X"06",X"36",X"36",X"33",X"C9",X"01",X"06",X"36",X"36",X"35",X"90",X"34",X"10",X"10",X"DF",X"77",
		X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"06",X"1F",X"03",X"20",X"89",X"34",X"10",X"CB",
		X"06",X"1F",X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"20",X"C2",X"34",X"10",X"10",
		X"DF",X"77",X"24",X"02",X"31",X"22",X"10",X"EE",X"22",X"CB",X"06",X"1F",X"03",X"7E",X"D2",X"AE",
		X"34",X"10",X"CB",X"06",X"1F",X"03",X"CC",X"00",X"00",X"8E",X"00",X"00",X"31",X"84",X"20",X"99",
		X"34",X"76",X"1A",X"01",X"09",X"8A",X"44",X"34",X"02",X"86",X"00",X"24",X"08",X"58",X"49",X"58",
		X"49",X"58",X"49",X"58",X"49",X"BD",X"D6",X"FE",X"DD",X"73",X"C6",X"03",X"E0",X"E0",X"A6",X"85",
		X"9B",X"74",X"19",X"A7",X"85",X"5A",X"2B",X"0E",X"A6",X"85",X"99",X"73",X"19",X"A7",X"85",X"86",
		X"00",X"97",X"73",X"5A",X"2A",X"F2",X"DC",X"AB",X"27",X"2B",X"30",X"01",X"31",X"03",X"8D",X"2A",
		X"25",X"23",X"A6",X"21",X"9B",X"AC",X"19",X"A7",X"21",X"A6",X"A4",X"99",X"AB",X"19",X"A7",X"A4",
		X"6C",X"06",X"6C",X"08",X"BD",X"D6",X"29",X"BD",X"D6",X"80",X"CC",X"D4",X"B0",X"BD",X"D5",X"4D",
		X"C6",X"05",X"BD",X"F5",X"1C",X"8D",X"12",X"35",X"76",X"39",X"34",X"06",X"EC",X"84",X"10",X"A3",
		X"A4",X"26",X"04",X"A6",X"02",X"A1",X"22",X"35",X"86",X"96",X"8B",X"34",X"02",X"4A",X"26",X"08",
		X"8E",X"0F",X"1C",X"CE",X"A1",X"C3",X"20",X"06",X"8E",X"71",X"1C",X"CE",X"A2",X"00",X"0F",X"73",
		X"C6",X"06",X"96",X"36",X"34",X"02",X"86",X"02",X"97",X"36",X"B7",X"D0",X"00",X"A6",X"C0",X"10",
		X"BE",X"C0",X"00",X"C5",X"01",X"26",X"06",X"33",X"5F",X"44",X"44",X"44",X"44",X"84",X"0F",X"26",
		X"0F",X"C1",X"02",X"23",X"0B",X"0D",X"73",X"26",X"07",X"1E",X"10",X"BD",X"F5",X"7B",X"20",X"0B",
		X"0C",X"73",X"48",X"48",X"31",X"A6",X"1E",X"10",X"BD",X"F5",X"22",X"1E",X"10",X"30",X"89",X"04",
		X"00",X"5A",X"26",X"C9",X"35",X"02",X"97",X"36",X"B7",X"D0",X"00",X"35",X"82",X"96",X"BA",X"2A",
		X"2A",X"BD",X"F5",X"07",X"BD",X"C0",X"33",X"7C",X"A1",X"62",X"20",X"1F",X"96",X"BA",X"2A",X"1B",
		X"1A",X"90",X"7F",X"D0",X"00",X"86",X"04",X"B7",X"CC",X"03",X"B6",X"CC",X"02",X"BD",X"F5",X"07",
		X"96",X"79",X"44",X"25",X"03",X"7E",X"C0",X"27",X"7E",X"C0",X"21",X"7E",X"D0",X"0A",X"8E",X"A0",
		X"7F",X"C6",X"12",X"20",X"0C",X"8E",X"A0",X"80",X"C6",X"15",X"20",X"05",X"8E",X"A0",X"81",X"C6",
		X"18",X"96",X"7E",X"26",X"E6",X"A6",X"84",X"26",X"E2",X"86",X"16",X"A7",X"84",X"86",X"C0",X"ED",
		X"49",X"86",X"0A",X"8E",X"D4",X"99",X"7E",X"D0",X"01",X"96",X"7E",X"26",X"CE",X"CC",X"D4",X"AB",
		X"BD",X"D5",X"4D",X"BD",X"F5",X"07",X"AD",X"D8",X"09",X"20",X"C0",X"FF",X"01",X"18",X"19",X"00",
		X"FF",X"01",X"20",X"1E",X"00",X"F0",X"02",X"08",X"11",X"01",X"20",X"17",X"00",X"F0",X"01",X"40",
		X"0A",X"00",X"F0",X"01",X"10",X"0B",X"00",X"E8",X"01",X"04",X"14",X"02",X"06",X"11",X"02",X"0A",
		X"17",X"00",X"E8",X"06",X"04",X"11",X"01",X"10",X"17",X"00",X"E0",X"03",X"0A",X"08",X"00",X"E0",
		X"01",X"18",X"1F",X"00",X"E0",X"01",X"18",X"11",X"00",X"D8",X"01",X"10",X"1A",X"00",X"D0",X"01",
		X"30",X"15",X"00",X"D0",X"01",X"10",X"05",X"00",X"D0",X"01",X"08",X"17",X"00",X"D0",X"01",X"08",
		X"07",X"00",X"D0",X"01",X"0A",X"01",X"00",X"D0",X"01",X"0A",X"06",X"00",X"D0",X"01",X"10",X"0B",
		X"00",X"C8",X"0A",X"01",X"0E",X"00",X"C0",X"01",X"08",X"07",X"00",X"C0",X"01",X"30",X"14",X"00",
		X"C0",X"01",X"20",X"18",X"00",X"C0",X"01",X"08",X"03",X"00",X"C0",X"01",X"30",X"09",X"00",X"C0",
		X"01",X"08",X"03",X"00",X"C0",X"01",X"18",X"0C",X"00",X"34",X"07",X"1A",X"FF",X"7F",X"D0",X"00",
		X"86",X"3F",X"B7",X"CC",X"02",X"53",X"C4",X"3F",X"F7",X"CC",X"02",X"35",X"87",X"34",X"17",X"0F",
		X"AD",X"1F",X"01",X"A6",X"84",X"91",X"B2",X"25",X"0D",X"97",X"B2",X"30",X"1E",X"1A",X"10",X"9F",
		X"B0",X"CC",X"01",X"01",X"DD",X"B3",X"35",X"97",X"96",X"B3",X"27",X"14",X"0A",X"B3",X"26",X"38",
		X"9E",X"B0",X"0A",X"B4",X"26",X"2C",X"30",X"03",X"9F",X"B0",X"A6",X"84",X"26",X"22",X"97",X"B2",
		X"96",X"7B",X"85",X"02",X"26",X"0A",X"96",X"AD",X"27",X"1E",X"0F",X"AD",X"C6",X"0F",X"20",X"16",
		X"96",X"AD",X"26",X"14",X"96",X"BA",X"85",X"98",X"26",X"0E",X"C6",X"16",X"D7",X"AD",X"20",X"06",
		X"97",X"B4",X"EC",X"01",X"97",X"B3",X"8D",X"91",X"B6",X"CC",X"01",X"85",X"40",X"27",X"04",X"86",
		X"3C",X"97",X"7E",X"96",X"7E",X"27",X"02",X"0A",X"7E",X"96",X"7F",X"27",X"02",X"0A",X"7F",X"96",
		X"81",X"27",X"02",X"0A",X"81",X"96",X"80",X"27",X"02",X"0A",X"80",X"96",X"7B",X"9A",X"7C",X"43",
		X"D6",X"7B",X"D7",X"7C",X"F6",X"CC",X"04",X"D7",X"7B",X"F6",X"CC",X"06",X"D7",X"7D",X"94",X"7B",
		X"27",X"1B",X"CE",X"F8",X"82",X"5F",X"CB",X"04",X"44",X"24",X"FB",X"33",X"C5",X"37",X"16",X"DE",
		X"82",X"26",X"05",X"DD",X"82",X"9F",X"84",X"39",X"DD",X"86",X"9F",X"88",X"39",X"96",X"79",X"9A",
		X"7A",X"43",X"D6",X"79",X"D7",X"7A",X"F6",X"CC",X"00",X"C4",X"3F",X"D7",X"79",X"95",X"79",X"27",
		X"17",X"8E",X"00",X"78",X"30",X"1F",X"26",X"FC",X"F6",X"CC",X"00",X"D4",X"79",X"D7",X"79",X"94",
		X"79",X"27",X"05",X"CE",X"F8",X"A2",X"8D",X"BD",X"39",X"34",X"76",X"8E",X"0F",X"14",X"B6",X"A1",
		X"C9",X"8D",X"0F",X"96",X"8C",X"4A",X"27",X"08",X"8E",X"71",X"14",X"B6",X"A2",X"06",X"8D",X"02",
		X"35",X"F6",X"81",X"05",X"23",X"02",X"86",X"05",X"34",X"02",X"CC",X"20",X"06",X"BD",X"F5",X"C7",
		X"A6",X"E4",X"27",X"0F",X"10",X"8E",X"F9",X"D5",X"1F",X"10",X"BD",X"F5",X"22",X"8B",X"06",X"6A",
		X"E4",X"26",X"F7",X"35",X"82",X"34",X"76",X"CC",X"40",X"20",X"8E",X"30",X"08",X"BD",X"F5",X"C7",
		X"8D",X"4A",X"8D",X"B5",X"8D",X"0A",X"96",X"8C",X"BD",X"D3",X"DB",X"4A",X"26",X"FA",X"35",X"F6",
		X"34",X"76",X"8E",X"29",X"1B",X"B6",X"A1",X"CB",X"8D",X"0F",X"96",X"8C",X"4A",X"27",X"08",X"8E",
		X"8B",X"1B",X"B6",X"A2",X"08",X"8D",X"02",X"35",X"F6",X"81",X"03",X"23",X"02",X"86",X"03",X"34",
		X"02",X"CC",X"03",X"0B",X"BD",X"F5",X"C7",X"A6",X"E4",X"27",X"0F",X"10",X"8E",X"F9",X"D9",X"1F",
		X"10",X"BD",X"F5",X"22",X"CB",X"04",X"6A",X"E4",X"26",X"F7",X"35",X"82",X"CC",X"55",X"55",X"8E",
		X"00",X"28",X"ED",X"84",X"30",X"89",X"01",X"00",X"8C",X"9C",X"00",X"25",X"F5",X"8E",X"2F",X"08",
		X"ED",X"89",X"41",X"00",X"ED",X"81",X"8C",X"2F",X"28",X"26",X"F5",X"8E",X"2F",X"07",X"A7",X"84",
		X"30",X"89",X"01",X"00",X"8C",X"71",X"07",X"26",X"F5",X"8E",X"4C",X"07",X"CC",X"99",X"99",X"ED",
		X"84",X"ED",X"88",X"21",X"30",X"89",X"01",X"00",X"8C",X"54",X"07",X"26",X"F2",X"39",X"34",X"02",
		X"96",X"8B",X"8E",X"A1",X"C2",X"4A",X"27",X"03",X"8E",X"A1",X"FF",X"35",X"82",X"34",X"02",X"20",
		X"F1",X"34",X"04",X"D6",X"DF",X"86",X"03",X"3D",X"CB",X"11",X"96",X"E1",X"44",X"44",X"44",X"98",
		X"E1",X"44",X"06",X"E0",X"06",X"E1",X"DB",X"E1",X"D9",X"E0",X"D7",X"DF",X"96",X"DF",X"35",X"84",
		X"C0",X"FF",X"00",X"00",X"14",X"05",X"34",X"3E",X"1A",X"FF",X"10",X"CE",X"BF",X"FF",X"86",X"A0",
		X"1F",X"8B",X"7F",X"D0",X"00",X"C6",X"04",X"CE",X"CC",X"00",X"8E",X"D7",X"30",X"6F",X"41",X"A6",
		X"80",X"A7",X"C1",X"A6",X"03",X"A7",X"5F",X"5A",X"26",X"F3",X"BD",X"F5",X"D1",X"8E",X"9C",X"00",
		X"6F",X"80",X"C6",X"38",X"F7",X"C3",X"FC",X"8C",X"C0",X"00",X"26",X"F4",X"7F",X"CC",X"00",X"7F",
		X"CC",X"02",X"8E",X"C4",X"7D",X"BD",X"F8",X"3A",X"1F",X"98",X"81",X"20",X"22",X"06",X"84",X"0F",
		X"81",X"09",X"23",X"01",X"5F",X"D7",X"37",X"CC",X"A5",X"5A",X"DD",X"E0",X"CC",X"FF",X"70",X"DD",
		X"A1",X"0F",X"A3",X"C6",X"FF",X"DD",X"79",X"BD",X"D8",X"DC",X"BD",X"F5",X"07",X"BD",X"C0",X"33",
		X"8D",X"24",X"8D",X"12",X"BD",X"F8",X"00",X"8E",X"D8",X"25",X"86",X"01",X"BD",X"D0",X"55",X"03",
		X"BA",X"1C",X"00",X"7E",X"E7",X"BE",X"8D",X"3D",X"BD",X"E6",X"9F",X"BD",X"E0",X"52",X"8D",X"45",
		X"BD",X"E5",X"4B",X"7E",X"E1",X"49",X"34",X"16",X"4F",X"5F",X"8E",X"AA",X"C5",X"9F",X"61",X"30",
		X"0F",X"AF",X"11",X"8C",X"AF",X"1B",X"26",X"F7",X"ED",X"84",X"DD",X"5F",X"8E",X"AF",X"2A",X"9F",
		X"69",X"30",X"88",X"17",X"AF",X"88",X"E9",X"8C",X"AF",X"86",X"26",X"F5",X"ED",X"84",X"8E",X"A0",
		X"5F",X"9F",X"63",X"35",X"96",X"8E",X"F8",X"BE",X"CE",X"A0",X"26",X"C6",X"10",X"A6",X"80",X"A7",
		X"C0",X"5A",X"26",X"F9",X"39",X"34",X"17",X"1A",X"FF",X"8E",X"A2",X"3C",X"9F",X"67",X"30",X"88",
		X"17",X"AF",X"88",X"E9",X"8C",X"AA",X"AE",X"26",X"F5",X"4F",X"5F",X"ED",X"84",X"DD",X"6B",X"DD",
		X"65",X"DD",X"6D",X"35",X"97",X"BD",X"F5",X"0B",X"7E",X"C0",X"00",X"8E",X"C4",X"95",X"BD",X"F8",
		X"22",X"4A",X"26",X"04",X"86",X"02",X"97",X"37",X"39",X"96",X"BA",X"2A",X"0E",X"8D",X"EC",X"96",
		X"37",X"27",X"08",X"CC",X"D4",X"BD",X"BD",X"D5",X"4D",X"8D",X"16",X"7E",X"D0",X"0A",X"96",X"BA",
		X"2A",X"F9",X"8D",X"D7",X"96",X"37",X"81",X"02",X"25",X"F1",X"8D",X"05",X"CC",X"D4",X"C2",X"20",
		X"E5",X"0F",X"38",X"12",X"96",X"B7",X"27",X"73",X"96",X"BA",X"2A",X"58",X"BD",X"D0",X"7C",X"BD",
		X"F5",X"D1",X"86",X"7F",X"97",X"BA",X"86",X"01",X"97",X"8B",X"97",X"25",X"0F",X"8C",X"8E",X"A1",
		X"C2",X"6F",X"80",X"8C",X"A2",X"3C",X"26",X"F9",X"8E",X"C4",X"85",X"BD",X"F8",X"22",X"84",X"0F",
		X"B7",X"A1",X"C9",X"C6",X"0A",X"FD",X"A1",X"CB",X"0F",X"39",X"12",X"8E",X"A1",X"C2",X"BD",X"DE",
		X"7C",X"8E",X"C4",X"81",X"BD",X"F8",X"38",X"DD",X"AB",X"FD",X"A1",X"C6",X"7F",X"A1",X"C8",X"8E",
		X"A1",X"C2",X"A6",X"80",X"A7",X"88",X"3C",X"8C",X"A1",X"FF",X"26",X"F6",X"8E",X"D9",X"19",X"86",
		X"00",X"BD",X"D0",X"55",X"0C",X"8C",X"96",X"37",X"8B",X"99",X"19",X"97",X"37",X"8E",X"C4",X"7D",
		X"BD",X"F8",X"4E",X"96",X"8C",X"4A",X"27",X"03",X"BD",X"D6",X"65",X"39",X"34",X"12",X"96",X"36",
		X"34",X"02",X"8E",X"DF",X"17",X"CC",X"38",X"3C",X"20",X"15",X"34",X"12",X"96",X"36",X"34",X"02",
		X"4F",X"BD",X"F5",X"0D",X"B6",X"CC",X"06",X"2A",X"E9",X"8E",X"DF",X"C3",X"CC",X"39",X"34",X"9F",
		X"90",X"0F",X"36",X"7F",X"D0",X"00",X"F7",X"CC",X"07",X"B7",X"C3",X"FC",X"86",X"7E",X"97",X"8F",
		X"35",X"02",X"97",X"36",X"B7",X"D0",X"00",X"35",X"92",X"C6",X"07",X"BD",X"F5",X"1C",X"BD",X"D7",
		X"B6",X"BD",X"D0",X"7C",X"86",X"7F",X"97",X"BA",X"9E",X"63",X"9C",X"5F",X"26",X"04",X"AE",X"84",
		X"27",X"10",X"86",X"0F",X"8E",X"D9",X"3A",X"7E",X"D0",X"01",X"96",X"7F",X"9A",X"80",X"9A",X"7F",
		X"26",X"F0",X"BD",X"D7",X"C6",X"8E",X"D9",X"50",X"86",X"00",X"BD",X"D0",X"55",X"7E",X"E7",X"BE",
		X"4F",X"BD",X"F5",X"0D",X"B6",X"CC",X"06",X"2A",X"15",X"BD",X"F5",X"D1",X"96",X"8B",X"4A",X"26",
		X"05",X"BD",X"D8",X"DC",X"20",X"02",X"8D",X"82",X"86",X"FF",X"97",X"7B",X"97",X"7C",X"4F",X"5F",
		X"DD",X"20",X"DD",X"22",X"BD",X"F4",X"FF",X"BD",X"C0",X"06",X"BD",X"C0",X"00",X"BD",X"F5",X"F1",
		X"CC",X"03",X"00",X"DD",X"BD",X"DD",X"BB",X"0F",X"AD",X"0F",X"B5",X"0F",X"8A",X"0F",X"AF",X"0F",
		X"9A",X"0F",X"99",X"8E",X"A1",X"1A",X"9F",X"9B",X"BD",X"D6",X"FE",X"9F",X"8D",X"A6",X"08",X"84",
		X"07",X"CE",X"DB",X"53",X"A6",X"C6",X"97",X"2B",X"6A",X"07",X"BD",X"D6",X"65",X"CC",X"20",X"80",
		X"DD",X"C1",X"DD",X"BF",X"CC",X"20",X"00",X"DD",X"C3",X"CC",X"08",X"00",X"D3",X"20",X"DD",X"CC",
		X"CC",X"80",X"00",X"DD",X"C5",X"4F",X"5F",X"DD",X"C7",X"97",X"C9",X"DD",X"CA",X"8E",X"E9",X"E3",
		X"86",X"00",X"BD",X"D0",X"55",X"8E",X"E7",X"82",X"86",X"00",X"BD",X"D0",X"55",X"8E",X"F4",X"93",
		X"86",X"00",X"BD",X"D0",X"55",X"8E",X"E9",X"BF",X"86",X"00",X"BD",X"D0",X"55",X"8E",X"F4",X"64",
		X"86",X"00",X"BD",X"D0",X"55",X"8E",X"F4",X"3D",X"86",X"00",X"BD",X"D0",X"55",X"96",X"25",X"27",
		X"1E",X"D6",X"8C",X"5A",X"27",X"19",X"CE",X"C0",X"EF",X"96",X"8B",X"4A",X"27",X"03",X"CE",X"C0",
		X"F1",X"8E",X"3C",X"80",X"BD",X"F5",X"13",X"86",X"80",X"8E",X"DA",X"1F",X"7E",X"D0",X"01",X"BD",
		X"F5",X"F1",X"C6",X"05",X"9E",X"8D",X"A6",X"0A",X"8D",X"15",X"86",X"60",X"8E",X"DA",X"32",X"7E",
		X"D0",X"01",X"BD",X"DC",X"1E",X"8D",X"05",X"0F",X"25",X"7E",X"DC",X"D9",X"5F",X"96",X"FA",X"26",
		X"02",X"CA",X"02",X"D7",X"BA",X"39",X"C6",X"58",X"8D",X"F3",X"DC",X"20",X"DD",X"22",X"9E",X"BF",
		X"CC",X"08",X"06",X"BD",X"F5",X"C7",X"BD",X"DB",X"B6",X"CC",X"D4",X"B5",X"BD",X"D5",X"4D",X"10",
		X"8E",X"F9",X"C1",X"96",X"BB",X"2A",X"04",X"10",X"8E",X"F9",X"CB",X"8E",X"DB",X"4B",X"AF",X"47",
		X"CE",X"AF",X"DD",X"BD",X"DB",X"5C",X"1F",X"31",X"DE",X"63",X"AF",X"4B",X"DC",X"C1",X"10",X"AE",
		X"4B",X"BD",X"F5",X"7B",X"86",X"02",X"8E",X"DA",X"8C",X"7E",X"D0",X"01",X"DC",X"C1",X"10",X"AE",
		X"4B",X"BD",X"F5",X"22",X"AE",X"47",X"A6",X"80",X"27",X"0E",X"97",X"31",X"0F",X"26",X"AF",X"47",
		X"86",X"02",X"8E",X"DA",X"7C",X"7E",X"D0",X"01",X"86",X"7F",X"97",X"BA",X"86",X"FF",X"97",X"26",
		X"86",X"02",X"8E",X"DA",X"B8",X"7E",X"D0",X"01",X"0F",X"26",X"BD",X"D0",X"7C",X"9E",X"C1",X"30",
		X"89",X"04",X"03",X"BD",X"F4",X"FF",X"BD",X"C0",X"0E",X"BD",X"D3",X"D9",X"0F",X"B3",X"C6",X"13",
		X"BD",X"D5",X"39",X"BD",X"DD",X"AE",X"26",X"06",X"BD",X"DD",X"EC",X"BD",X"F5",X"F1",X"96",X"8B",
		X"9E",X"8D",X"E6",X"07",X"26",X"2F",X"D6",X"8C",X"5A",X"27",X"41",X"88",X"03",X"BD",X"D7",X"0D",
		X"E6",X"07",X"27",X"38",X"CE",X"C0",X"EF",X"81",X"02",X"27",X"03",X"CE",X"C0",X"F1",X"8E",X"3C",
		X"78",X"BD",X"F5",X"13",X"CE",X"C0",X"75",X"8E",X"3E",X"88",X"BD",X"F5",X"13",X"86",X"60",X"8E",
		X"DB",X"15",X"7E",X"D0",X"01",X"96",X"8B",X"4C",X"91",X"8C",X"23",X"02",X"86",X"01",X"BD",X"D7",
		X"0D",X"E6",X"07",X"27",X"F2",X"97",X"8B",X"0C",X"25",X"7E",X"D9",X"19",X"CE",X"C0",X"75",X"8E",
		X"3E",X"80",X"86",X"FF",X"97",X"BA",X"BD",X"F5",X"13",X"0F",X"B3",X"C6",X"13",X"BD",X"D5",X"39",
		X"86",X"28",X"8E",X"DB",X"48",X"7E",X"D0",X"01",X"7E",X"D8",X"25",X"07",X"07",X"07",X"0F",X"3F",
		X"7F",X"FF",X"FF",X"00",X"81",X"28",X"07",X"16",X"2F",X"84",X"15",X"00",X"34",X"56",X"BD",X"F5",
		X"03",X"EC",X"A4",X"ED",X"C4",X"3D",X"30",X"4A",X"AF",X"42",X"30",X"8B",X"AF",X"44",X"34",X"10",
		X"30",X"8B",X"34",X"10",X"EC",X"26",X"ED",X"46",X"EC",X"28",X"ED",X"48",X"AE",X"22",X"33",X"4A",
		X"8D",X"0E",X"AE",X"24",X"EE",X"62",X"EC",X"E4",X"ED",X"62",X"8D",X"04",X"32",X"64",X"35",X"D6",
		X"EC",X"81",X"85",X"F0",X"27",X"02",X"8A",X"F0",X"85",X"0F",X"27",X"02",X"8A",X"0F",X"C5",X"F0",
		X"27",X"02",X"CA",X"F0",X"C5",X"0F",X"27",X"02",X"CA",X"0F",X"84",X"BB",X"C4",X"BB",X"ED",X"C1",
		X"11",X"A3",X"64",X"25",X"DB",X"39",X"34",X"56",X"DE",X"8D",X"33",X"4A",X"86",X"33",X"6F",X"C0",
		X"4A",X"26",X"FB",X"DE",X"8D",X"96",X"FA",X"A7",X"4A",X"33",X"4B",X"8E",X"A0",X"FB",X"A6",X"80",
		X"8C",X"A1",X"00",X"22",X"03",X"AB",X"88",X"16",X"A7",X"C0",X"8C",X"A1",X"12",X"26",X"EF",X"35",
		X"D6",X"34",X"06",X"97",X"74",X"BD",X"D0",X"95",X"F9",X"01",X"ED",X"70",X"66",X"66",X"BD",X"D7",
		X"11",X"DC",X"E0",X"84",X"1F",X"AB",X"61",X"ED",X"0A",X"54",X"24",X"05",X"CC",X"F9",X"15",X"ED",
		X"02",X"86",X"E0",X"A7",X"0C",X"86",X"10",X"A7",X"88",X"14",X"4F",X"5F",X"ED",X"88",X"10",X"ED",
		X"0E",X"ED",X"06",X"9F",X"65",X"AF",X"A1",X"0A",X"74",X"26",X"CA",X"35",X"86",X"0C",X"8E",X"EC",
		X"C9",X"86",X"00",X"BD",X"D0",X"55",X"CE",X"A1",X"1A",X"31",X"C4",X"EF",X"07",X"6F",X"C0",X"11",
		X"83",X"A1",X"42",X"26",X"F8",X"DE",X"8D",X"A6",X"4A",X"97",X"FA",X"27",X"20",X"81",X"07",X"23",
		X"10",X"44",X"44",X"5F",X"8D",X"9B",X"CB",X"40",X"26",X"FA",X"48",X"48",X"40",X"AB",X"4A",X"27",
		X"0C",X"97",X"73",X"D6",X"E0",X"86",X"01",X"8D",X"88",X"0A",X"73",X"26",X"F6",X"DE",X"8D",X"33",
		X"4B",X"8E",X"A0",X"FB",X"A6",X"C0",X"A7",X"80",X"8C",X"A1",X"12",X"26",X"F7",X"8E",X"A1",X"12",
		X"6F",X"80",X"8C",X"A1",X"1A",X"26",X"F9",X"BD",X"D0",X"AD",X"96",X"DF",X"44",X"8B",X"2A",X"A7",
		X"0C",X"BD",X"D7",X"11",X"84",X"3F",X"8B",X"80",X"D3",X"20",X"ED",X"0A",X"96",X"FF",X"27",X"19",
		X"81",X"06",X"23",X"02",X"86",X"06",X"31",X"84",X"BD",X"EB",X"9E",X"9E",X"67",X"AF",X"A4",X"10",
		X"9F",X"67",X"40",X"9B",X"FF",X"97",X"FF",X"26",X"CE",X"96",X"FE",X"27",X"05",X"BD",X"EF",X"15",
		X"0F",X"FE",X"96",X"FD",X"B7",X"A1",X"14",X"27",X"05",X"0F",X"FD",X"BD",X"EB",X"36",X"96",X"FC",
		X"B7",X"A1",X"13",X"27",X"13",X"81",X"03",X"23",X"02",X"86",X"03",X"34",X"02",X"BD",X"F2",X"9D",
		X"96",X"FC",X"A0",X"E0",X"97",X"FC",X"26",X"ED",X"39",X"DE",X"63",X"86",X"28",X"A7",X"47",X"B6",
		X"A1",X"0F",X"B7",X"A1",X"18",X"86",X"01",X"B7",X"A1",X"17",X"96",X"BA",X"85",X"08",X"26",X"7C",
		X"BD",X"DD",X"AE",X"26",X"14",X"86",X"77",X"97",X"BA",X"BD",X"D0",X"7C",X"BD",X"DB",X"B6",X"BD",
		X"DD",X"EC",X"9E",X"8D",X"6C",X"07",X"7E",X"D9",X"1E",X"81",X"08",X"22",X"12",X"F6",X"A1",X"0F",
		X"54",X"81",X"03",X"22",X"01",X"54",X"5C",X"F1",X"A1",X"18",X"24",X"03",X"F7",X"A1",X"18",X"7A",
		X"A1",X"18",X"26",X"1C",X"81",X"04",X"B6",X"A1",X"0F",X"24",X"05",X"44",X"44",X"BD",X"DD",X"9E",
		X"B7",X"A1",X"18",X"B6",X"A1",X"19",X"81",X"0C",X"24",X"06",X"BD",X"EA",X"80",X"7C",X"A1",X"19",
		X"7A",X"A1",X"17",X"27",X"05",X"B6",X"A1",X"12",X"26",X"22",X"B6",X"A1",X"00",X"B7",X"A1",X"17",
		X"96",X"FB",X"27",X"18",X"B6",X"A1",X"12",X"81",X"08",X"24",X"11",X"B6",X"A1",X"01",X"91",X"FB",
		X"23",X"02",X"96",X"FB",X"BD",X"EF",X"9C",X"40",X"9B",X"FB",X"97",X"FB",X"96",X"AE",X"81",X"10",
		X"24",X"02",X"0C",X"AE",X"96",X"24",X"4C",X"81",X"F0",X"23",X"06",X"C6",X"06",X"BD",X"F5",X"1C",
		X"4F",X"97",X"24",X"DE",X"63",X"6A",X"47",X"26",X"0D",X"C6",X"02",X"10",X"8E",X"A0",X"FB",X"BD",
		X"DE",X"EC",X"86",X"28",X"A7",X"47",X"86",X"0F",X"8E",X"DC",X"EA",X"7E",X"D0",X"01",X"34",X"02",
		X"BD",X"D7",X"11",X"A1",X"E4",X"23",X"03",X"44",X"20",X"F9",X"4C",X"32",X"61",X"39",X"B6",X"A1",
		X"12",X"9B",X"FB",X"BB",X"A1",X"13",X"BB",X"A1",X"14",X"BB",X"A1",X"16",X"BB",X"A1",X"15",X"9B",
		X"FE",X"39",X"34",X"04",X"5F",X"81",X"10",X"25",X"06",X"CB",X"0A",X"80",X"10",X"20",X"F6",X"34",
		X"04",X"AB",X"E0",X"35",X"84",X"34",X"04",X"1F",X"89",X"4F",X"C1",X"0A",X"25",X"07",X"8B",X"10",
		X"19",X"C0",X"0A",X"20",X"F5",X"34",X"04",X"AB",X"E0",X"19",X"35",X"84",X"0F",X"26",X"DE",X"63",
		X"35",X"10",X"AF",X"4D",X"BD",X"F5",X"F1",X"CE",X"C0",X"F9",X"8E",X"38",X"50",X"BD",X"F5",X"13",
		X"9E",X"8D",X"A6",X"08",X"8D",X"CF",X"1F",X"89",X"4F",X"9E",X"50",X"BD",X"C0",X"0E",X"8E",X"3D",
		X"60",X"CE",X"C0",X"FB",X"BD",X"F5",X"13",X"CE",X"C0",X"F3",X"8E",X"3C",X"90",X"BD",X"F5",X"13",
		X"9E",X"8D",X"5F",X"A6",X"08",X"81",X"05",X"23",X"02",X"86",X"05",X"9E",X"50",X"BD",X"C0",X"0E",
		X"DE",X"63",X"8E",X"3C",X"A0",X"96",X"FA",X"A7",X"49",X"27",X"31",X"1F",X"10",X"10",X"8E",X"F9",
		X"15",X"BD",X"F5",X"22",X"30",X"89",X"04",X"00",X"86",X"01",X"10",X"9E",X"8D",X"E6",X"28",X"C1",
		X"05",X"25",X"02",X"C6",X"05",X"58",X"58",X"58",X"58",X"BD",X"D3",X"60",X"AF",X"47",X"86",X"04",
		X"8E",X"DE",X"66",X"7E",X"D0",X"01",X"AE",X"47",X"6A",X"49",X"26",X"CF",X"9E",X"8D",X"BD",X"DE",
		X"7C",X"86",X"80",X"8E",X"DE",X"79",X"7E",X"D0",X"01",X"6E",X"D8",X"0D",X"34",X"56",X"6C",X"08",
		X"8E",X"C4",X"9D",X"BD",X"F8",X"22",X"97",X"73",X"AE",X"62",X"4D",X"27",X"0C",X"A6",X"08",X"90",
		X"73",X"25",X"06",X"26",X"FA",X"86",X"0A",X"A7",X"0A",X"BD",X"F4",X"FF",X"A6",X"08",X"34",X"02",
		X"81",X"04",X"23",X"02",X"86",X"04",X"FE",X"C0",X"11",X"8B",X"03",X"30",X"0B",X"E6",X"C6",X"E7",
		X"80",X"33",X"48",X"11",X"B3",X"C0",X"13",X"26",X"F4",X"35",X"02",X"80",X"04",X"24",X"01",X"4F",
		X"97",X"73",X"8E",X"C4",X"97",X"BD",X"F8",X"38",X"BD",X"DD",X"C2",X"9B",X"73",X"97",X"73",X"27",
		X"19",X"1F",X"98",X"BD",X"DD",X"C2",X"91",X"73",X"24",X"02",X"97",X"73",X"96",X"73",X"C6",X"03",
		X"BD",X"D6",X"FE",X"31",X"0B",X"8D",X"05",X"4A",X"26",X"F4",X"35",X"D6",X"34",X"32",X"BD",X"F4",
		X"FF",X"BE",X"C0",X"11",X"A6",X"85",X"2B",X"0A",X"AB",X"A4",X"25",X"10",X"A1",X"84",X"22",X"0C",
		X"20",X"08",X"AB",X"A4",X"24",X"06",X"A1",X"01",X"25",X"02",X"A7",X"A4",X"31",X"21",X"30",X"08",
		X"BC",X"C0",X"13",X"26",X"DF",X"35",X"B2",X"7F",X"D0",X"00",X"86",X"A0",X"1F",X"8B",X"86",X"04",
		X"B7",X"CC",X"03",X"B6",X"CC",X"02",X"B6",X"C8",X"00",X"81",X"80",X"25",X"30",X"96",X"92",X"26",
		X"7B",X"0C",X"92",X"BD",X"D5",X"68",X"BD",X"E2",X"63",X"BD",X"E0",X"7E",X"B6",X"C8",X"00",X"80",
		X"08",X"81",X"A8",X"23",X"02",X"86",X"A8",X"97",X"A2",X"86",X"02",X"B7",X"D0",X"00",X"DC",X"A2",
		X"BD",X"E3",X"9F",X"DC",X"A2",X"BD",X"E2",X"13",X"BD",X"E4",X"53",X"20",X"4F",X"D6",X"92",X"27",
		X"4B",X"0F",X"92",X"0C",X"5D",X"C6",X"38",X"F7",X"C3",X"FC",X"81",X"08",X"22",X"1B",X"CE",X"C0",
		X"10",X"DC",X"30",X"9E",X"32",X"10",X"9E",X"34",X"36",X"36",X"DC",X"2A",X"9E",X"2C",X"10",X"9E",
		X"2E",X"36",X"36",X"DC",X"26",X"9E",X"28",X"36",X"16",X"BD",X"D5",X"FD",X"86",X"07",X"B7",X"D0",
		X"00",X"96",X"BA",X"85",X"02",X"26",X"03",X"BD",X"C0",X"03",X"86",X"02",X"B7",X"D0",X"00",X"DC",
		X"A1",X"BD",X"E2",X"13",X"DC",X"A1",X"BD",X"E3",X"9F",X"BD",X"E3",X"76",X"1A",X"FF",X"7F",X"D0",
		X"00",X"86",X"05",X"B7",X"CC",X"03",X"96",X"36",X"B7",X"D0",X"00",X"A6",X"E4",X"84",X"6F",X"A7",
		X"E4",X"35",X"FF",X"7F",X"D0",X"00",X"86",X"A0",X"1F",X"8B",X"86",X"04",X"B7",X"CC",X"03",X"B6",
		X"CC",X"02",X"B6",X"C8",X"00",X"81",X"58",X"25",X"2C",X"D6",X"92",X"26",X"CF",X"0C",X"92",X"43",
		X"12",X"97",X"A2",X"BD",X"D5",X"FD",X"86",X"07",X"B7",X"D0",X"00",X"96",X"BA",X"85",X"02",X"26",
		X"03",X"BD",X"C0",X"03",X"86",X"02",X"B7",X"D0",X"00",X"DC",X"A1",X"BD",X"E2",X"13",X"DC",X"A1",
		X"BD",X"E3",X"9F",X"20",X"A7",X"D6",X"92",X"27",X"A3",X"0F",X"92",X"0C",X"5D",X"C6",X"39",X"F7",
		X"C3",X"FC",X"81",X"04",X"22",X"1B",X"CE",X"C0",X"10",X"DC",X"30",X"9E",X"32",X"10",X"9E",X"34",
		X"36",X"36",X"DC",X"2A",X"9E",X"2C",X"10",X"9E",X"2E",X"36",X"36",X"DC",X"26",X"9E",X"28",X"36",
		X"16",X"BD",X"D5",X"68",X"BD",X"E2",X"63",X"BD",X"E0",X"7E",X"86",X"02",X"B7",X"D0",X"00",X"DC",
		X"A2",X"BD",X"E2",X"13",X"DC",X"A2",X"BD",X"E3",X"9F",X"BD",X"E4",X"53",X"BD",X"E3",X"76",X"7E",
		X"DF",X"AC",X"8E",X"AF",X"9D",X"C6",X"10",X"D7",X"AE",X"5F",X"BD",X"D7",X"11",X"81",X"9C",X"24",
		X"F9",X"A7",X"84",X"BD",X"D7",X"11",X"81",X"A8",X"22",X"F9",X"81",X"2A",X"23",X"F5",X"A7",X"01",
		X"E7",X"02",X"CB",X"11",X"C4",X"77",X"30",X"04",X"8C",X"AF",X"DD",X"26",X"DD",X"39",X"96",X"BA",
		X"85",X"20",X"26",X"F9",X"8E",X"AF",X"9D",X"DC",X"20",X"C4",X"80",X"DD",X"6F",X"DC",X"22",X"C4",
		X"80",X"93",X"6F",X"58",X"49",X"97",X"6F",X"C6",X"F0",X"96",X"21",X"85",X"40",X"26",X"01",X"53",
		X"D7",X"71",X"4F",X"A7",X"94",X"A7",X"98",X"04",X"A7",X"98",X"08",X"A7",X"98",X"0C",X"A7",X"98",
		X"10",X"A7",X"98",X"14",X"A7",X"98",X"18",X"A7",X"98",X"1C",X"A7",X"98",X"20",X"A7",X"98",X"24",
		X"A7",X"98",X"28",X"A7",X"98",X"2C",X"A7",X"98",X"30",X"A7",X"98",X"34",X"A7",X"98",X"38",X"A7",
		X"98",X"3C",X"D6",X"AE",X"A6",X"84",X"9B",X"6F",X"81",X"9C",X"25",X"0A",X"81",X"C0",X"23",X"04",
		X"86",X"9B",X"20",X"02",X"86",X"00",X"A7",X"84",X"A6",X"02",X"94",X"71",X"A7",X"98",X"00",X"30",
		X"04",X"5A",X"26",X"E0",X"D6",X"DF",X"C4",X"3C",X"8E",X"AF",X"9D",X"3A",X"A6",X"02",X"8B",X"11",
		X"84",X"77",X"A7",X"02",X"96",X"DF",X"85",X"01",X"26",X"3E",X"81",X"98",X"25",X"24",X"CE",X"A1",
		X"02",X"33",X"C8",X"B6",X"EE",X"C4",X"11",X"83",X"62",X"45",X"27",X"14",X"0D",X"BA",X"2B",X"10",
		X"81",X"A0",X"25",X"0C",X"81",X"A1",X"24",X"08",X"D6",X"E1",X"1F",X"01",X"D6",X"E0",X"E7",X"84",
		X"80",X"84",X"6F",X"98",X"00",X"A7",X"84",X"96",X"BA",X"85",X"02",X"27",X"0B",X"96",X"E1",X"84",
		X"3F",X"C6",X"03",X"3D",X"CB",X"2A",X"E7",X"01",X"39",X"8E",X"A1",X"62",X"9F",X"9F",X"BD",X"D7",
		X"11",X"A7",X"88",X"20",X"A7",X"80",X"8C",X"A1",X"83",X"26",X"F3",X"39",X"9E",X"9F",X"DE",X"BF",
		X"33",X"C9",X"FF",X"01",X"EC",X"84",X"ED",X"C4",X"A6",X"05",X"E6",X"09",X"ED",X"42",X"A6",X"0C",
		X"A7",X"44",X"96",X"7B",X"85",X"02",X"27",X"22",X"A6",X"03",X"E6",X"06",X"ED",X"C9",X"FF",X"01",
		X"A6",X"0A",X"A7",X"C9",X"FF",X"03",X"A6",X"04",X"E6",X"07",X"ED",X"C9",X"FE",X"01",X"A6",X"0B",
		X"A7",X"C9",X"FE",X"03",X"A6",X"08",X"A7",X"C9",X"FD",X"02",X"39",X"DE",X"9F",X"9E",X"BF",X"30",
		X"89",X"08",X"01",X"37",X"26",X"ED",X"84",X"10",X"AF",X"02",X"37",X"26",X"A7",X"04",X"96",X"7B",
		X"85",X"02",X"27",X"18",X"E7",X"89",X"01",X"01",X"10",X"AF",X"89",X"01",X"02",X"37",X"26",X"10",
		X"AF",X"89",X"02",X"01",X"A7",X"89",X"02",X"03",X"E7",X"89",X"03",X"02",X"39",X"DE",X"BF",X"5F",
		X"8E",X"00",X"00",X"31",X"84",X"33",X"C9",X"08",X"06",X"36",X"34",X"AF",X"C9",X"01",X"01",X"E7",
		X"C9",X"01",X"03",X"AF",X"C9",X"02",X"01",X"E7",X"C9",X"02",X"03",X"E7",X"C9",X"03",X"02",X"39",
		X"DE",X"BF",X"5F",X"8E",X"00",X"00",X"31",X"84",X"33",X"C9",X"FF",X"06",X"36",X"34",X"AF",X"C9",
		X"FF",X"01",X"E7",X"C9",X"FF",X"03",X"AF",X"C9",X"FE",X"01",X"E7",X"C9",X"FE",X"03",X"E7",X"C9",
		X"FD",X"02",X"39",X"97",X"77",X"96",X"BA",X"85",X"10",X"26",X"28",X"96",X"77",X"91",X"C0",X"23",
		X"22",X"D1",X"C0",X"22",X"1E",X"96",X"BD",X"2B",X"08",X"BD",X"E2",X"5E",X"BD",X"E1",X"F0",X"20",
		X"06",X"BD",X"E2",X"5E",X"BD",X"E1",X"CD",X"DC",X"BB",X"DD",X"BD",X"2B",X"07",X"BD",X"E2",X"4A",
		X"BD",X"E1",X"5C",X"39",X"BD",X"E2",X"58",X"7E",X"E1",X"9B",X"10",X"8E",X"F9",X"C1",X"96",X"C4",
		X"48",X"DC",X"C1",X"DD",X"BF",X"7E",X"D2",X"8E",X"10",X"8E",X"F9",X"CB",X"20",X"F0",X"DC",X"BF",
		X"7E",X"D2",X"DF",X"96",X"BA",X"85",X"40",X"10",X"26",X"01",X"0A",X"0F",X"6F",X"DC",X"C7",X"43",
		X"53",X"C3",X"00",X"01",X"2A",X"02",X"03",X"6F",X"58",X"49",X"58",X"49",X"D3",X"C8",X"DD",X"C8",
		X"96",X"6F",X"99",X"C7",X"97",X"C7",X"DC",X"C7",X"96",X"7B",X"85",X"02",X"27",X"12",X"0F",X"6F",
		X"DC",X"BD",X"2A",X"02",X"03",X"6F",X"D3",X"C8",X"DD",X"C8",X"96",X"6F",X"99",X"C7",X"97",X"C7",
		X"DC",X"C7",X"47",X"56",X"47",X"56",X"4F",X"57",X"46",X"97",X"94",X"D7",X"93",X"96",X"BD",X"2B",
		X"07",X"86",X"20",X"5D",X"2B",X"07",X"20",X"09",X"86",X"70",X"5D",X"2B",X"04",X"0F",X"94",X"0F",
		X"93",X"D6",X"94",X"9B",X"93",X"97",X"93",X"93",X"C3",X"27",X"26",X"25",X"12",X"10",X"83",X"01",
		X"00",X"23",X"1E",X"CC",X"00",X"40",X"DD",X"95",X"CC",X"01",X"00",X"D3",X"C3",X"20",X"18",X"10",
		X"83",X"FF",X"00",X"2E",X"0C",X"CC",X"FF",X"C0",X"DD",X"95",X"CC",X"FF",X"00",X"D3",X"C3",X"20",
		X"06",X"4F",X"5F",X"DD",X"95",X"DC",X"93",X"DD",X"C3",X"97",X"C1",X"DC",X"20",X"DD",X"22",X"DC",
		X"C7",X"10",X"83",X"01",X"00",X"2D",X"03",X"CC",X"01",X"00",X"10",X"83",X"FF",X"00",X"2E",X"03",
		X"CC",X"FF",X"00",X"DD",X"C7",X"D3",X"20",X"93",X"95",X"DD",X"20",X"DC",X"C3",X"44",X"56",X"44",
		X"56",X"C4",X"E0",X"D3",X"20",X"DD",X"CC",X"D6",X"C5",X"96",X"7D",X"44",X"25",X"09",X"96",X"7B",
		X"2B",X"20",X"CC",X"00",X"00",X"20",X"36",X"C1",X"2B",X"23",X"3A",X"DC",X"CA",X"2A",X"0E",X"C3",
		X"FF",X"F8",X"10",X"83",X"FE",X"00",X"2C",X"25",X"CC",X"FE",X"00",X"20",X"20",X"CC",X"FF",X"00",
		X"20",X"1B",X"C1",X"EE",X"24",X"1F",X"DC",X"CA",X"2F",X"0E",X"C3",X"00",X"08",X"10",X"83",X"02",
		X"00",X"23",X"0A",X"CC",X"02",X"00",X"20",X"05",X"CC",X"01",X"00",X"20",X"00",X"DD",X"CA",X"D3",
		X"C5",X"DD",X"C5",X"97",X"C2",X"39",X"96",X"BA",X"85",X"20",X"26",X"22",X"8E",X"A0",X"65",X"20",
		X"19",X"EC",X"0A",X"E3",X"0E",X"ED",X"0A",X"EC",X"0C",X"E3",X"88",X"10",X"81",X"2A",X"24",X"02",
		X"86",X"F0",X"81",X"F0",X"23",X"02",X"86",X"2A",X"ED",X"0C",X"AE",X"84",X"26",X"E3",X"39",X"34",
		X"06",X"96",X"BA",X"85",X"20",X"26",X"4A",X"8E",X"A0",X"65",X"20",X"41",X"EC",X"04",X"27",X"12",
		X"E1",X"E4",X"22",X"39",X"E1",X"61",X"23",X"35",X"10",X"AE",X"02",X"AD",X"B8",X"08",X"4F",X"5F",
		X"ED",X"04",X"E6",X"0C",X"E1",X"E4",X"22",X"25",X"E1",X"61",X"23",X"21",X"EC",X"0A",X"93",X"20",
		X"10",X"83",X"25",X"80",X"24",X"17",X"10",X"AE",X"02",X"58",X"49",X"58",X"49",X"AB",X"A4",X"81",
		X"9C",X"22",X"0A",X"A0",X"A4",X"58",X"E6",X"0C",X"ED",X"04",X"AD",X"B8",X"06",X"AE",X"84",X"26",
		X"BB",X"35",X"86",X"34",X"66",X"96",X"99",X"81",X"14",X"24",X"4F",X"EC",X"0A",X"93",X"20",X"10",
		X"83",X"25",X"80",X"24",X"45",X"58",X"49",X"58",X"49",X"E6",X"0C",X"C1",X"2A",X"23",X"3B",X"9E",
		X"67",X"27",X"37",X"ED",X"04",X"ED",X"0A",X"1E",X"89",X"ED",X"0C",X"EF",X"06",X"4F",X"5F",X"ED",
		X"0E",X"ED",X"88",X"10",X"EE",X"66",X"37",X"26",X"ED",X"88",X"12",X"10",X"AF",X"02",X"37",X"06",
		X"EF",X"66",X"ED",X"08",X"86",X"14",X"A7",X"88",X"15",X"A7",X"88",X"16",X"EC",X"84",X"DD",X"67",
		X"DC",X"6D",X"ED",X"84",X"0C",X"99",X"9F",X"6D",X"35",X"E6",X"EE",X"66",X"33",X"46",X"EF",X"66",
		X"4F",X"35",X"E6",X"96",X"BA",X"85",X"20",X"26",X"3E",X"DC",X"20",X"C4",X"E0",X"DD",X"9D",X"DC",
		X"22",X"C4",X"E0",X"93",X"9D",X"58",X"49",X"58",X"49",X"DD",X"9D",X"8E",X"A0",X"6D",X"20",X"23",
		X"10",X"AE",X"04",X"EC",X"88",X"10",X"E3",X"0C",X"81",X"2A",X"23",X"4A",X"ED",X"0C",X"EC",X"0E",
		X"D3",X"9D",X"E3",X"0A",X"81",X"98",X"24",X"3E",X"ED",X"0A",X"E6",X"0C",X"ED",X"04",X"EE",X"04",
		X"6E",X"98",X"12",X"AE",X"84",X"26",X"D9",X"39",X"DE",X"A6",X"E6",X"0B",X"2A",X"02",X"33",X"46",
		X"CC",X"00",X"00",X"ED",X"A4",X"A7",X"22",X"ED",X"A9",X"01",X"00",X"A7",X"A9",X"01",X"02",X"10",
		X"AE",X"04",X"EC",X"C4",X"ED",X"A4",X"EC",X"42",X"A7",X"22",X"E7",X"A9",X"01",X"00",X"EC",X"44",
		X"ED",X"A9",X"01",X"01",X"20",X"CD",X"4F",X"5F",X"A7",X"88",X"16",X"ED",X"A4",X"A7",X"22",X"ED",
		X"A9",X"01",X"00",X"A7",X"A9",X"01",X"02",X"20",X"BA",X"DE",X"A8",X"E6",X"0B",X"58",X"CC",X"00",
		X"00",X"ED",X"A4",X"A7",X"22",X"ED",X"A9",X"01",X"00",X"A7",X"A9",X"01",X"02",X"10",X"AE",X"04",
		X"25",X"15",X"EC",X"C4",X"84",X"0F",X"ED",X"A4",X"EC",X"42",X"84",X"0F",X"A7",X"22",X"C4",X"F0",
		X"E7",X"A9",X"01",X"01",X"7E",X"E4",X"93",X"EC",X"C4",X"C4",X"0F",X"E7",X"21",X"84",X"F0",X"A7",
		X"A9",X"01",X"02",X"EC",X"42",X"84",X"F0",X"ED",X"A9",X"01",X"00",X"7E",X"E4",X"93",X"CC",X"00",
		X"25",X"BD",X"D3",X"60",X"0A",X"99",X"BD",X"D0",X"F2",X"BD",X"F3",X"FE",X"EC",X"0A",X"44",X"56",
		X"44",X"56",X"D3",X"20",X"ED",X"0A",X"A6",X"0C",X"80",X"02",X"A7",X"0C",X"CC",X"F9",X"51",X"ED",
		X"02",X"BD",X"FC",X"63",X"CC",X"D4",X"E4",X"7E",X"D5",X"4D",X"5E",X"8E",X"A1",X"A2",X"9F",X"A8",
		X"C6",X"0A",X"BD",X"D7",X"11",X"2B",X"02",X"C6",X"09",X"44",X"25",X"04",X"CB",X"A0",X"20",X"02",
		X"CB",X"90",X"E7",X"80",X"8C",X"A1",X"C2",X"26",X"E7",X"39",X"8E",X"A0",X"6D",X"20",X"1B",X"A6",
		X"88",X"16",X"27",X"05",X"6A",X"88",X"15",X"26",X"11",X"EE",X"84",X"EF",X"A4",X"DE",X"67",X"EF",
		X"84",X"9F",X"67",X"BD",X"F3",X"FE",X"0A",X"99",X"30",X"A4",X"31",X"84",X"AE",X"84",X"26",X"DF",
		X"39",X"96",X"B5",X"81",X"04",X"24",X"11",X"0C",X"B5",X"CC",X"D5",X"1B",X"BD",X"D5",X"4D",X"9E",
		X"C1",X"96",X"BB",X"2A",X"1C",X"7E",X"E6",X"30",X"7E",X"D0",X"0A",X"34",X"46",X"86",X"02",X"97",
		X"36",X"B7",X"D0",X"00",X"35",X"06",X"12",X"12",X"12",X"CE",X"F9",X"6F",X"BD",X"E6",X"BA",X"35",
		X"C0",X"30",X"89",X"07",X"04",X"AF",X"47",X"AF",X"49",X"AF",X"4B",X"96",X"BA",X"85",X"40",X"26",
		X"50",X"86",X"04",X"AE",X"47",X"C6",X"11",X"8C",X"98",X"00",X"24",X"45",X"E7",X"84",X"30",X"89",
		X"01",X"00",X"4A",X"26",X"F7",X"C6",X"99",X"E7",X"84",X"AF",X"47",X"10",X"9E",X"A4",X"10",X"8C",
		X"A1",X"5F",X"25",X"04",X"10",X"8E",X"A1",X"42",X"AE",X"49",X"86",X"03",X"E6",X"A0",X"E7",X"84",
		X"30",X"89",X"01",X"00",X"4A",X"26",X"F5",X"10",X"9F",X"A4",X"AF",X"49",X"6F",X"D8",X"0B",X"6C",
		X"4B",X"EC",X"47",X"80",X"06",X"8D",X"94",X"26",X"08",X"86",X"01",X"8E",X"E5",X"CB",X"7E",X"D0",
		X"01",X"AE",X"4B",X"4F",X"A7",X"84",X"30",X"89",X"01",X"00",X"AC",X"47",X"23",X"F6",X"20",X"6A",
		X"30",X"04",X"AF",X"47",X"AF",X"49",X"AF",X"4B",X"96",X"BA",X"85",X"40",X"26",X"4F",X"86",X"04",
		X"AE",X"47",X"C6",X"11",X"8C",X"05",X"00",X"23",X"44",X"E7",X"84",X"30",X"89",X"FF",X"00",X"4A",
		X"26",X"F7",X"C6",X"99",X"E7",X"84",X"AF",X"47",X"10",X"9E",X"A4",X"10",X"8C",X"A1",X"5F",X"25",
		X"04",X"10",X"8E",X"A1",X"42",X"AE",X"49",X"86",X"03",X"E6",X"A0",X"E7",X"84",X"30",X"89",X"FF",
		X"00",X"4A",X"26",X"F5",X"10",X"9F",X"A4",X"AF",X"49",X"6F",X"D8",X"0B",X"6A",X"4B",X"EC",X"47",
		X"BD",X"E5",X"AB",X"26",X"08",X"86",X"01",X"8E",X"E6",X"38",X"7E",X"D0",X"01",X"AE",X"4B",X"4F",
		X"A7",X"84",X"30",X"89",X"FF",X"00",X"AC",X"47",X"24",X"F6",X"0A",X"B5",X"7E",X"D0",X"0A",X"8E",
		X"A1",X"42",X"9F",X"A4",X"BD",X"D7",X"11",X"5F",X"44",X"24",X"02",X"CB",X"01",X"44",X"24",X"02",
		X"CB",X"10",X"E7",X"80",X"8C",X"A1",X"62",X"26",X"EB",X"39",X"8E",X"A0",X"65",X"DD",X"D6",X"E3",
		X"C4",X"DD",X"D8",X"20",X"17",X"EC",X"04",X"27",X"13",X"91",X"D8",X"24",X"0F",X"D1",X"D9",X"24",
		X"0B",X"E3",X"98",X"02",X"91",X"D6",X"23",X"04",X"D1",X"D7",X"22",X"05",X"AE",X"84",X"26",X"E5",
		X"39",X"DF",X"DC",X"10",X"AE",X"02",X"A3",X"A4",X"DD",X"73",X"4F",X"5F",X"DD",X"D0",X"DD",X"D2",
		X"DC",X"73",X"D0",X"D7",X"22",X"05",X"50",X"D7",X"D1",X"20",X"02",X"D7",X"D3",X"90",X"D6",X"22",
		X"05",X"40",X"97",X"D0",X"20",X"02",X"97",X"D2",X"DC",X"73",X"E3",X"A4",X"D0",X"D9",X"22",X"01",
		X"5F",X"90",X"D8",X"22",X"01",X"4F",X"DD",X"DA",X"EC",X"A4",X"93",X"D0",X"93",X"DA",X"DD",X"CE",
		X"A6",X"41",X"97",X"D5",X"D6",X"D2",X"3D",X"EE",X"42",X"33",X"CB",X"A6",X"21",X"97",X"D4",X"10",
		X"AE",X"22",X"D6",X"D0",X"3D",X"31",X"AB",X"96",X"D1",X"31",X"A6",X"96",X"D3",X"33",X"C6",X"D6",
		X"CF",X"5A",X"A6",X"C5",X"27",X"2A",X"A6",X"A5",X"27",X"26",X"31",X"A5",X"1F",X"20",X"EE",X"02",
		X"A3",X"42",X"10",X"AE",X"04",X"E0",X"41",X"82",X"00",X"25",X"06",X"31",X"A9",X"01",X"00",X"20",
		X"F4",X"EB",X"41",X"89",X"00",X"31",X"A5",X"10",X"9F",X"F8",X"AD",X"98",X"08",X"86",X"01",X"39",
		X"5A",X"2A",X"CF",X"DC",X"D4",X"31",X"A6",X"33",X"C5",X"0A",X"CE",X"26",X"C2",X"DE",X"DC",X"7E",
		X"E6",X"DC",X"0F",X"B6",X"8E",X"E7",X"99",X"96",X"B6",X"E6",X"86",X"27",X"F5",X"0C",X"B6",X"D7",
		X"27",X"86",X"02",X"8E",X"E7",X"84",X"7E",X"D0",X"01",X"38",X"39",X"3A",X"3B",X"3C",X"3D",X"3E",
		X"3F",X"37",X"2F",X"27",X"1F",X"17",X"47",X"47",X"87",X"87",X"C7",X"C7",X"C6",X"C5",X"CC",X"CB",
		X"CA",X"DA",X"E8",X"F8",X"F9",X"FA",X"FB",X"FD",X"FF",X"BF",X"3F",X"3E",X"3C",X"00",X"8E",X"A0",
		X"5F",X"9F",X"63",X"96",X"5D",X"27",X"FC",X"0F",X"5D",X"D6",X"BA",X"C5",X"7D",X"27",X"04",X"0F",
		X"5E",X"20",X"47",X"48",X"9B",X"5E",X"80",X"04",X"2A",X"01",X"4F",X"97",X"5E",X"81",X"02",X"25",
		X"39",X"C6",X"03",X"D7",X"AE",X"81",X"02",X"23",X"31",X"86",X"02",X"97",X"5E",X"10",X"8E",X"A0",
		X"65",X"AE",X"A4",X"27",X"25",X"A6",X"88",X"14",X"27",X"04",X"31",X"84",X"20",X"F3",X"EE",X"84",
		X"EF",X"A4",X"DC",X"DF",X"84",X"3F",X"8B",X"60",X"E3",X"0A",X"ED",X"0A",X"BD",X"F3",X"FE",X"CC",
		X"00",X"00",X"ED",X"04",X"DE",X"6B",X"9F",X"6B",X"EF",X"84",X"86",X"02",X"97",X"36",X"B7",X"D0",
		X"00",X"8D",X"3E",X"BD",X"FC",X"66",X"BD",X"D7",X"11",X"9E",X"82",X"26",X"0C",X"9E",X"86",X"27",
		X"17",X"DC",X"88",X"0F",X"86",X"0F",X"87",X"20",X"06",X"DC",X"84",X"0F",X"82",X"0F",X"83",X"D4",
		X"BA",X"26",X"E6",X"BD",X"D0",X"55",X"20",X"E1",X"CE",X"A0",X"5F",X"20",X"09",X"6A",X"44",X"26",
		X"05",X"DF",X"63",X"6E",X"D8",X"02",X"EE",X"C4",X"26",X"F3",X"10",X"CE",X"BF",X"FF",X"7E",X"E7",
		X"BE",X"96",X"BA",X"85",X"10",X"26",X"2D",X"DC",X"BF",X"CE",X"F9",X"C1",X"0D",X"BD",X"2A",X"03",
		X"CE",X"F9",X"CB",X"34",X"46",X"0C",X"DE",X"BD",X"E6",X"BA",X"35",X"46",X"26",X"08",X"8E",X"A0",
		X"6D",X"BD",X"E6",X"BD",X"27",X"0E",X"8E",X"DA",X"46",X"86",X"00",X"BD",X"D0",X"55",X"96",X"BA",
		X"8A",X"08",X"97",X"BA",X"0F",X"DE",X"39",X"96",X"AF",X"26",X"23",X"0C",X"AF",X"DC",X"BD",X"53",
		X"43",X"C3",X"00",X"01",X"DD",X"BB",X"86",X"02",X"8E",X"E8",X"AE",X"7E",X"D0",X"01",X"96",X"7B",
		X"85",X"40",X"26",X"F2",X"86",X"05",X"8E",X"E8",X"BC",X"7E",X"D0",X"01",X"0F",X"AF",X"7E",X"D0",
		X"0A",X"96",X"9A",X"26",X"57",X"9E",X"8D",X"A6",X"09",X"27",X"51",X"0C",X"9A",X"6A",X"09",X"BD",
		X"D6",X"80",X"CC",X"D4",X"D2",X"BD",X"D5",X"4D",X"9E",X"65",X"27",X"14",X"EC",X"04",X"27",X"0C",
		X"A6",X"88",X"14",X"81",X"02",X"24",X"05",X"AD",X"98",X"08",X"20",X"EC",X"AE",X"84",X"20",X"EA",
		X"DE",X"63",X"86",X"04",X"A7",X"47",X"03",X"26",X"86",X"02",X"8E",X"E9",X"00",X"7E",X"D0",X"01",
		X"6A",X"47",X"26",X"F2",X"86",X"0A",X"8E",X"E9",X"0C",X"7E",X"D0",X"01",X"96",X"7B",X"85",X"04",
		X"26",X"F2",X"86",X"0A",X"8E",X"E9",X"1A",X"7E",X"D0",X"01",X"0F",X"9A",X"7E",X"D0",X"0A",X"96",
		X"BA",X"85",X"FD",X"10",X"26",X"00",X"95",X"86",X"77",X"97",X"BA",X"BD",X"F5",X"F1",X"86",X"0F",
		X"8E",X"E9",X"36",X"7E",X"D0",X"01",X"9E",X"6D",X"27",X"05",X"BD",X"D0",X"F2",X"20",X"F7",X"0F",
		X"99",X"DC",X"DF",X"DD",X"20",X"DD",X"22",X"54",X"24",X"08",X"CC",X"20",X"00",X"8E",X"03",X"00",
		X"20",X"06",X"8E",X"FD",X"00",X"CC",X"70",X"00",X"DD",X"C3",X"9F",X"BB",X"D6",X"E0",X"54",X"CB",
		X"2A",X"D7",X"C5",X"DD",X"C1",X"4F",X"5F",X"97",X"C9",X"DD",X"C7",X"DD",X"CA",X"BD",X"F4",X"FA",
		X"C6",X"50",X"BD",X"DA",X"3D",X"BD",X"D0",X"95",X"F9",X"C1",X"ED",X"BC",X"00",X"00",X"CC",X"00",
		X"00",X"ED",X"0E",X"ED",X"88",X"10",X"DC",X"C5",X"ED",X"0C",X"DC",X"C3",X"44",X"56",X"44",X"56",
		X"D3",X"20",X"ED",X"0A",X"96",X"BB",X"2A",X"05",X"CE",X"F9",X"CB",X"EF",X"02",X"DE",X"63",X"AF",
		X"47",X"BD",X"FC",X"60",X"86",X"28",X"8E",X"E9",X"AC",X"7E",X"D0",X"01",X"AE",X"47",X"BD",X"F3",
		X"FB",X"BD",X"DA",X"3C",X"96",X"E1",X"81",X"C0",X"10",X"22",X"F0",X"8A",X"7E",X"D0",X"0A",X"9E",
		X"9F",X"30",X"01",X"8C",X"A1",X"82",X"23",X"03",X"8E",X"A1",X"62",X"9F",X"9F",X"9E",X"A8",X"30",
		X"01",X"8C",X"A1",X"BA",X"23",X"03",X"8E",X"A1",X"A2",X"9F",X"A8",X"86",X"04",X"8E",X"E9",X"BF",
		X"7E",X"D0",X"01",X"BD",X"EA",X"33",X"86",X"02",X"8E",X"E9",X"EE",X"7E",X"D0",X"01",X"BD",X"EA",
		X"0A",X"BD",X"E5",X"6A",X"86",X"02",X"8E",X"E9",X"FC",X"7E",X"D0",X"01",X"BD",X"F5",X"0B",X"BD",
		X"C0",X"03",X"86",X"04",X"8E",X"E9",X"E3",X"7E",X"D0",X"01",X"DC",X"20",X"83",X"0C",X"80",X"DD",
		X"73",X"8E",X"A0",X"65",X"20",X"16",X"EC",X"0A",X"93",X"73",X"10",X"83",X"3E",X"80",X"25",X"0C",
		X"EE",X"84",X"EF",X"A4",X"DE",X"6B",X"EF",X"84",X"9F",X"6B",X"30",X"A4",X"31",X"84",X"AE",X"84",
		X"26",X"E4",X"39",X"DC",X"20",X"83",X"0C",X"80",X"DD",X"73",X"8E",X"A0",X"6B",X"20",X"39",X"EC",
		X"88",X"10",X"58",X"49",X"58",X"49",X"58",X"49",X"E3",X"0C",X"81",X"2A",X"24",X"02",X"86",X"F0",
		X"81",X"F0",X"23",X"02",X"86",X"2A",X"ED",X"0C",X"EC",X"0E",X"58",X"49",X"58",X"49",X"58",X"49",
		X"E3",X"0A",X"ED",X"0A",X"93",X"73",X"10",X"83",X"3E",X"80",X"24",X"0C",X"EE",X"84",X"EF",X"A4",
		X"DE",X"65",X"EF",X"84",X"9F",X"65",X"30",X"A4",X"31",X"84",X"AE",X"84",X"26",X"C1",X"39",X"40",
		X"8E",X"EA",X"B4",X"86",X"00",X"BD",X"D0",X"55",X"33",X"84",X"BD",X"D0",X"95",X"F9",X"A3",X"EB",
		X"2B",X"33",X"33",X"AF",X"47",X"EF",X"06",X"DC",X"DF",X"84",X"1F",X"D3",X"20",X"ED",X"0A",X"54",
		X"CB",X"2A",X"E7",X"0C",X"4F",X"5F",X"ED",X"88",X"10",X"ED",X"0E",X"86",X"08",X"A7",X"49",X"8D",
		X"44",X"7E",X"FC",X"60",X"AE",X"47",X"EC",X"02",X"10",X"83",X"F8",X"EC",X"27",X"28",X"6A",X"49",
		X"26",X"13",X"B6",X"A1",X"10",X"BD",X"DD",X"9E",X"A7",X"49",X"BD",X"EE",X"BA",X"27",X"06",X"CC",
		X"D5",X"2F",X"BD",X"D5",X"4D",X"EE",X"02",X"33",X"4A",X"11",X"83",X"F9",X"B7",X"23",X"05",X"CE",
		X"F9",X"A3",X"8D",X"0A",X"EF",X"02",X"86",X"06",X"8E",X"EA",X"B4",X"7E",X"D0",X"01",X"96",X"DF",
		X"B1",X"A1",X"11",X"23",X"35",X"CC",X"40",X"01",X"DD",X"73",X"EC",X"0A",X"93",X"CC",X"2B",X"02",
		X"00",X"73",X"C3",X"02",X"80",X"10",X"83",X"05",X"00",X"23",X"07",X"D6",X"73",X"1D",X"D3",X"C7",
		X"ED",X"0E",X"A6",X"0C",X"90",X"C0",X"2B",X"02",X"00",X"74",X"8B",X"0A",X"81",X"14",X"23",X"0A",
		X"5F",X"96",X"74",X"D3",X"CA",X"47",X"56",X"ED",X"88",X"10",X"39",X"7A",X"A1",X"19",X"BD",X"F4",
		X"16",X"01",X"20",X"D4",X"FD",X"39",X"97",X"73",X"BD",X"D0",X"95",X"F8",X"F7",X"EB",X"74",X"CC",
		X"CC",X"BD",X"D7",X"11",X"DC",X"E0",X"84",X"3F",X"8B",X"10",X"ED",X"0A",X"54",X"CB",X"2A",X"E7",
		X"0C",X"D6",X"DF",X"C4",X"3F",X"CB",X"E0",X"1D",X"ED",X"0E",X"D6",X"E1",X"C4",X"7F",X"C0",X"40",
		X"1D",X"2B",X"04",X"CA",X"20",X"20",X"02",X"C4",X"DF",X"ED",X"88",X"10",X"BD",X"FC",X"60",X"0A",
		X"73",X"26",X"C5",X"39",X"BD",X"F4",X"1D",X"02",X"10",X"D4",X"F3",X"86",X"06",X"BD",X"DD",X"9E",
		X"31",X"84",X"BD",X"EB",X"9E",X"7A",X"A1",X"14",X"39",X"BD",X"D7",X"11",X"D6",X"DF",X"1D",X"58",
		X"49",X"ED",X"88",X"10",X"D6",X"E1",X"C4",X"3F",X"CB",X"E0",X"1D",X"ED",X"0E",X"39",X"34",X"76",
		X"97",X"73",X"B6",X"A1",X"16",X"4C",X"81",X"14",X"22",X"3D",X"B7",X"A1",X"16",X"8E",X"EC",X"17",
		X"86",X"00",X"BD",X"D0",X"55",X"33",X"84",X"BD",X"D0",X"95",X"F9",X"7B",X"EB",X"E9",X"24",X"24",
		X"EC",X"2A",X"ED",X"0A",X"EC",X"2C",X"ED",X"0C",X"AF",X"47",X"EF",X"06",X"8D",X"BB",X"DC",X"E0",
		X"F4",X"A1",X"0E",X"E7",X"49",X"84",X"1F",X"A7",X"44",X"B6",X"A1",X"0D",X"BD",X"DD",X"9E",X"A7",
		X"4B",X"9F",X"65",X"0A",X"73",X"26",X"BB",X"35",X"F6",X"7A",X"A1",X"16",X"BD",X"F3",X"FB",X"34",
		X"10",X"BD",X"D0",X"13",X"35",X"10",X"EC",X"0A",X"83",X"00",X"40",X"ED",X"0A",X"EC",X"0C",X"80",
		X"02",X"A7",X"0C",X"CE",X"F8",X"E2",X"EF",X"02",X"BD",X"FC",X"63",X"CC",X"01",X"15",X"BD",X"D3",
		X"60",X"CC",X"D5",X"16",X"7E",X"D5",X"4D",X"AE",X"47",X"F6",X"A1",X"0C",X"10",X"9E",X"CC",X"10",
		X"AC",X"0A",X"24",X"01",X"50",X"1D",X"ED",X"0E",X"20",X"54",X"E6",X"49",X"AE",X"47",X"96",X"C0",
		X"A1",X"0C",X"22",X"01",X"50",X"1D",X"E3",X"88",X"10",X"10",X"83",X"02",X"00",X"2D",X"03",X"CC",
		X"02",X"00",X"10",X"83",X"FE",X"00",X"2E",X"03",X"CC",X"FE",X"00",X"ED",X"88",X"10",X"43",X"53",
		X"58",X"49",X"58",X"49",X"1F",X"89",X"1D",X"E3",X"88",X"10",X"ED",X"88",X"10",X"D6",X"DF",X"C4",
		X"1F",X"CB",X"F0",X"1D",X"E3",X"88",X"10",X"ED",X"88",X"10",X"DC",X"CC",X"A3",X"0A",X"C3",X"12",
		X"C0",X"10",X"83",X"25",X"80",X"22",X"A0",X"6A",X"4B",X"26",X"03",X"BD",X"EC",X"86",X"86",X"03",
		X"8E",X"EC",X"2A",X"7E",X"D0",X"01",X"34",X"10",X"DC",X"CC",X"A3",X"0A",X"A8",X"0E",X"2B",X"2F",
		X"31",X"84",X"BD",X"E3",X"F3",X"E4",X"D9",X"F9",X"5B",X"E5",X"1E",X"27",X"22",X"EC",X"2E",X"58",
		X"49",X"58",X"49",X"58",X"49",X"ED",X"0E",X"CC",X"D5",X"34",X"BD",X"D5",X"4D",X"5F",X"96",X"C0",
		X"A0",X"0C",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"47",X"56",X"ED",X"88",X"10",X"B6",
		X"A1",X"0D",X"BD",X"DD",X"9E",X"A7",X"4B",X"35",X"90",X"AE",X"47",X"30",X"02",X"8C",X"A1",X"3A",
		X"25",X"03",X"8E",X"A1",X"1A",X"AF",X"47",X"AE",X"84",X"27",X"76",X"EC",X"04",X"27",X"72",X"EC",
		X"08",X"10",X"83",X"ED",X"70",X"26",X"6A",X"EC",X"02",X"10",X"83",X"F9",X"0B",X"22",X"2F",X"96",
		X"DF",X"81",X"08",X"23",X"50",X"BD",X"ED",X"59",X"8B",X"04",X"81",X"E8",X"23",X"02",X"86",X"E8",
		X"C6",X"01",X"A1",X"0C",X"27",X"07",X"22",X"01",X"50",X"EB",X"0C",X"E7",X"0C",X"EE",X"02",X"33",
		X"4A",X"11",X"83",X"F9",X"0B",X"23",X"03",X"CE",X"F9",X"01",X"C6",X"E0",X"20",X"2C",X"96",X"DF",
		X"81",X"08",X"23",X"F3",X"8D",X"33",X"8B",X"0F",X"81",X"E8",X"23",X"02",X"86",X"E8",X"C6",X"01",
		X"A1",X"0C",X"27",X"07",X"22",X"01",X"50",X"EB",X"0C",X"E7",X"0C",X"EE",X"02",X"33",X"4A",X"11",
		X"83",X"F9",X"1F",X"23",X"03",X"CE",X"F9",X"15",X"C6",X"20",X"EF",X"02",X"1D",X"E3",X"0A",X"ED",
		X"0A",X"86",X"02",X"8E",X"EC",X"C9",X"7E",X"D0",X"01",X"34",X"14",X"EC",X"0A",X"44",X"56",X"44",
		X"56",X"44",X"56",X"44",X"56",X"44",X"56",X"44",X"56",X"8E",X"B3",X"00",X"A6",X"8B",X"35",X"94",
		X"96",X"DE",X"27",X"03",X"4F",X"35",X"86",X"8D",X"4B",X"BD",X"F3",X"FB",X"CC",X"F8",X"D8",X"ED",
		X"02",X"EC",X"0A",X"83",X"00",X"40",X"ED",X"0A",X"BD",X"FC",X"63",X"CC",X"D4",X"E4",X"7E",X"D5",
		X"4D",X"EE",X"06",X"27",X"DB",X"96",X"DE",X"27",X"26",X"EC",X"42",X"10",X"83",X"F2",X"4C",X"27",
		X"16",X"CC",X"D4",X"DA",X"BD",X"D5",X"4D",X"34",X"10",X"8E",X"EE",X"73",X"86",X"00",X"BD",X"D0",
		X"55",X"31",X"84",X"35",X"10",X"AF",X"27",X"CC",X"F2",X"4C",X"ED",X"42",X"4F",X"35",X"86",X"8D",
		X"B6",X"7E",X"D0",X"13",X"31",X"84",X"34",X"52",X"CE",X"A1",X"1A",X"86",X"40",X"10",X"AC",X"C1",
		X"27",X"06",X"4A",X"26",X"F8",X"BD",X"D0",X"3A",X"4F",X"5F",X"ED",X"5E",X"0A",X"FA",X"26",X"08",
		X"8E",X"ED",X"EA",X"86",X"00",X"BD",X"D0",X"55",X"35",X"D2",X"96",X"BA",X"8A",X"02",X"97",X"BA",
		X"6F",X"47",X"BD",X"F4",X"FF",X"BD",X"C0",X"09",X"8E",X"B1",X"25",X"CE",X"00",X"00",X"86",X"40",
		X"EF",X"91",X"4A",X"26",X"FB",X"9E",X"67",X"CC",X"F9",X"F1",X"ED",X"02",X"C6",X"02",X"D7",X"73",
		X"BD",X"D7",X"11",X"84",X"3F",X"D3",X"20",X"ED",X"0A",X"BD",X"ED",X"59",X"A7",X"0C",X"80",X"0A",
		X"BD",X"FC",X"63",X"0A",X"73",X"26",X"E9",X"96",X"DF",X"84",X"1F",X"8E",X"E7",X"99",X"A6",X"86",
		X"97",X"26",X"CC",X"D4",X"E4",X"BD",X"D5",X"4D",X"8E",X"EE",X"44",X"86",X"02",X"C6",X"08",X"D7",
		X"5E",X"7E",X"D0",X"01",X"0F",X"26",X"A6",X"47",X"44",X"44",X"44",X"4C",X"BD",X"DD",X"9E",X"8E",
		X"EE",X"54",X"20",X"E9",X"6C",X"47",X"A6",X"47",X"81",X"10",X"26",X"A9",X"CC",X"D4",X"C7",X"BD",
		X"D5",X"4D",X"7E",X"D0",X"0A",X"BD",X"D0",X"95",X"F9",X"DD",X"ED",X"BC",X"00",X"00",X"CC",X"01",
		X"25",X"20",X"0C",X"BD",X"D0",X"95",X"F9",X"E7",X"ED",X"BC",X"00",X"00",X"CC",X"01",X"50",X"BD",
		X"D3",X"60",X"10",X"AE",X"47",X"DC",X"C7",X"ED",X"0E",X"CC",X"00",X"00",X"ED",X"88",X"10",X"86",
		X"11",X"A7",X"88",X"14",X"EC",X"2A",X"ED",X"0A",X"EC",X"2C",X"2B",X"05",X"C3",X"18",X"00",X"20",
		X"03",X"83",X"20",X"00",X"ED",X"0C",X"9F",X"65",X"AF",X"47",X"86",X"32",X"8E",X"EE",X"B2",X"7E",
		X"D0",X"01",X"AE",X"47",X"BD",X"F3",X"FB",X"7E",X"D0",X"0A",X"34",X"10",X"BD",X"E3",X"F3",X"E4",
		X"D9",X"F9",X"5B",X"E5",X"1E",X"27",X"35",X"D6",X"DF",X"C4",X"1F",X"CB",X"F0",X"DB",X"BF",X"E0",
		X"04",X"1D",X"58",X"49",X"58",X"49",X"ED",X"0E",X"D6",X"DF",X"C1",X"78",X"23",X"0A",X"DC",X"C7",
		X"58",X"49",X"58",X"49",X"E3",X"0E",X"ED",X"0E",X"D6",X"E1",X"C4",X"1F",X"CB",X"F0",X"DB",X"C0",
		X"E0",X"05",X"1D",X"58",X"49",X"58",X"49",X"ED",X"88",X"10",X"86",X"01",X"35",X"90",X"6A",X"4D",
		X"26",X"12",X"B6",X"A1",X"05",X"BD",X"DD",X"9E",X"A7",X"4D",X"8D",X"AE",X"27",X"06",X"CC",X"D5",
		X"25",X"BD",X"D5",X"4D",X"39",X"34",X"02",X"97",X"73",X"8E",X"F1",X"5E",X"86",X"00",X"BD",X"D0",
		X"55",X"33",X"84",X"BD",X"D0",X"95",X"F8",X"CE",X"EF",X"6D",X"CC",X"33",X"BD",X"D7",X"11",X"DC",
		X"20",X"83",X"25",X"80",X"DD",X"75",X"DC",X"E0",X"93",X"75",X"10",X"83",X"4B",X"00",X"24",X"03",
		X"C3",X"80",X"00",X"D3",X"75",X"ED",X"0A",X"96",X"DF",X"44",X"8B",X"2A",X"A7",X"0C",X"4F",X"5F",
		X"ED",X"88",X"10",X"ED",X"0E",X"B6",X"A1",X"0B",X"BD",X"DD",X"9E",X"A7",X"47",X"BD",X"FC",X"60",
		X"EF",X"06",X"AF",X"47",X"7C",X"A1",X"15",X"0A",X"73",X"26",X"AE",X"35",X"82",X"7A",X"A1",X"15",
		X"BD",X"F4",X"16",X"01",X"15",X"D4",X"F8",X"39",X"34",X"10",X"96",X"FA",X"27",X"1C",X"9E",X"9B",
		X"30",X"02",X"8C",X"A1",X"5A",X"25",X"03",X"8E",X"A1",X"1A",X"EC",X"84",X"26",X"06",X"9C",X"9B",
		X"26",X"EE",X"35",X"90",X"9F",X"9B",X"ED",X"49",X"AF",X"4B",X"35",X"90",X"34",X"02",X"97",X"73",
		X"0D",X"FA",X"26",X"03",X"7E",X"EF",X"19",X"8E",X"EF",X"F6",X"86",X"00",X"BD",X"D0",X"55",X"33",
		X"84",X"BD",X"D0",X"95",X"F9",X"85",X"F2",X"0B",X"44",X"33",X"BD",X"D7",X"11",X"DC",X"E0",X"ED",
		X"0A",X"86",X"2C",X"A7",X"0C",X"FC",X"A1",X"03",X"ED",X"88",X"10",X"B6",X"A1",X"05",X"BD",X"DD",
		X"9E",X"A7",X"4D",X"B6",X"A1",X"02",X"BD",X"DD",X"9E",X"1F",X"89",X"4F",X"C5",X"01",X"27",X"02",
		X"53",X"43",X"ED",X"0E",X"EF",X"06",X"BD",X"FC",X"60",X"AF",X"47",X"8D",X"8B",X"7C",X"A1",X"12",
		X"0A",X"73",X"26",X"AC",X"35",X"82",X"AE",X"47",X"10",X"AE",X"49",X"EC",X"D8",X"0B",X"27",X"16",
		X"A6",X"29",X"81",X"70",X"26",X"10",X"A6",X"0A",X"84",X"FC",X"97",X"73",X"A6",X"2A",X"84",X"FC",
		X"91",X"73",X"27",X"51",X"20",X"0F",X"A6",X"88",X"14",X"84",X"FE",X"A7",X"88",X"14",X"BD",X"EF",
		X"78",X"10",X"27",X"01",X"19",X"BD",X"ED",X"59",X"80",X"32",X"A0",X"0C",X"22",X"0F",X"81",X"EC",
		X"2D",X"04",X"4F",X"5F",X"20",X"0A",X"FC",X"A1",X"03",X"43",X"53",X"20",X"03",X"FC",X"A1",X"03",
		X"ED",X"88",X"10",X"EC",X"02",X"10",X"83",X"F8",X"EC",X"27",X"12",X"BD",X"EE",X"FE",X"EE",X"02",
		X"33",X"4A",X"11",X"83",X"F9",X"99",X"23",X"03",X"CE",X"F9",X"85",X"EF",X"02",X"86",X"06",X"8E",
		X"EF",X"F6",X"7E",X"D0",X"01",X"4F",X"5F",X"6C",X"88",X"14",X"ED",X"0E",X"ED",X"88",X"10",X"CC",
		X"F9",X"85",X"ED",X"02",X"AE",X"47",X"10",X"AE",X"49",X"EC",X"D8",X"0B",X"27",X"98",X"A6",X"29",
		X"81",X"70",X"26",X"92",X"EC",X"2A",X"C4",X"E0",X"DD",X"75",X"EC",X"0A",X"C4",X"E0",X"10",X"93",
		X"75",X"27",X"0D",X"2D",X"04",X"C6",X"E0",X"20",X"02",X"C6",X"20",X"1D",X"E3",X"0A",X"ED",X"0A",
		X"A6",X"2C",X"80",X"0C",X"A1",X"0C",X"27",X"16",X"FC",X"A1",X"03",X"24",X"02",X"43",X"53",X"E3",
		X"0C",X"ED",X"0C",X"BD",X"EE",X"FE",X"86",X"01",X"8E",X"F0",X"74",X"7E",X"D0",X"01",X"EC",X"0A",
		X"C3",X"00",X"40",X"A3",X"2A",X"10",X"83",X"00",X"80",X"22",X"E8",X"CC",X"F1",X"E0",X"ED",X"08",
		X"FC",X"A1",X"03",X"53",X"43",X"ED",X"88",X"10",X"ED",X"A8",X"10",X"CC",X"D5",X"0C",X"BD",X"D5",
		X"4D",X"CC",X"ED",X"91",X"ED",X"28",X"DE",X"63",X"AE",X"47",X"A6",X"0C",X"81",X"32",X"23",X"0B",
		X"BD",X"EE",X"FE",X"86",X"04",X"8E",X"F0",X"E6",X"7E",X"D0",X"01",X"CC",X"D5",X"11",X"BD",X"D5",
		X"4D",X"AE",X"47",X"10",X"AE",X"49",X"EC",X"D8",X"0B",X"26",X"0B",X"BD",X"F3",X"FB",X"7A",X"A1",
		X"12",X"0C",X"FB",X"7E",X"D0",X"0A",X"4F",X"5F",X"ED",X"88",X"10",X"ED",X"A8",X"10",X"A6",X"2C",
		X"A1",X"0C",X"23",X"0F",X"6A",X"2C",X"86",X"12",X"BD",X"D5",X"39",X"86",X"01",X"8E",X"F1",X"01",
		X"7E",X"D0",X"01",X"30",X"A4",X"EC",X"24",X"8B",X"01",X"DD",X"F8",X"BD",X"ED",X"77",X"7A",X"A1",
		X"12",X"7C",X"A1",X"15",X"AE",X"47",X"6F",X"88",X"14",X"CC",X"F8",X"CE",X"ED",X"02",X"CC",X"CC",
		X"33",X"ED",X"88",X"12",X"CC",X"EF",X"6D",X"ED",X"08",X"B6",X"A1",X"0B",X"A7",X"49",X"AE",X"47",
		X"F6",X"A1",X"0A",X"10",X"9E",X"CC",X"10",X"AC",X"0A",X"2C",X"01",X"50",X"1D",X"ED",X"0E",X"DC",
		X"CC",X"A3",X"0A",X"C3",X"01",X"7C",X"10",X"83",X"07",X"00",X"23",X"21",X"96",X"C0",X"A0",X"0C",
		X"23",X"0B",X"81",X"08",X"22",X"0B",X"FC",X"A1",X"08",X"43",X"53",X"20",X"0B",X"81",X"F8",X"2E",
		X"04",X"4F",X"5F",X"20",X"03",X"FC",X"A1",X"08",X"ED",X"88",X"10",X"20",X"12",X"96",X"C0",X"A1",
		X"0C",X"FC",X"A1",X"08",X"24",X"02",X"43",X"53",X"ED",X"88",X"10",X"EC",X"04",X"27",X"29",X"F6",
		X"A1",X"07",X"96",X"DF",X"2B",X"01",X"50",X"EB",X"0C",X"C1",X"2A",X"24",X"02",X"C6",X"F0",X"E7",
		X"0C",X"6A",X"49",X"26",X"13",X"B6",X"A1",X"0B",X"BD",X"DD",X"9E",X"A7",X"49",X"BD",X"EE",X"BA",
		X"27",X"06",X"CC",X"D5",X"2A",X"BD",X"D5",X"4D",X"86",X"03",X"8E",X"F1",X"5E",X"7E",X"D0",X"01",
		X"EE",X"06",X"EC",X"D8",X"0B",X"27",X"24",X"CC",X"00",X"00",X"CC",X"00",X"00",X"34",X"10",X"8E",
		X"F2",X"16",X"86",X"00",X"BD",X"D0",X"55",X"EE",X"49",X"EF",X"07",X"CC",X"D4",X"E9",X"BD",X"D5",
		X"4D",X"CC",X"00",X"00",X"ED",X"C8",X"10",X"AF",X"46",X"35",X"10",X"7A",X"A1",X"12",X"BD",X"F4",
		X"16",X"01",X"15",X"D5",X"07",X"39",X"AE",X"47",X"CC",X"00",X"08",X"E3",X"88",X"10",X"10",X"83",
		X"03",X"00",X"24",X"03",X"ED",X"88",X"10",X"BD",X"ED",X"59",X"A1",X"0C",X"22",X"16",X"EC",X"88",
		X"10",X"10",X"83",X"00",X"E0",X"23",X"39",X"EC",X"04",X"C3",X"01",X"07",X"DD",X"F8",X"BD",X"ED",
		X"77",X"7E",X"D0",X"0A",X"86",X"04",X"8E",X"F2",X"16",X"7E",X"D0",X"01",X"AE",X"47",X"CC",X"00",
		X"00",X"ED",X"88",X"10",X"96",X"C5",X"8B",X"0A",X"A7",X"0C",X"DC",X"CC",X"C3",X"00",X"80",X"ED",
		X"0A",X"BD",X"ED",X"59",X"A1",X"0C",X"25",X"0F",X"86",X"01",X"8E",X"F2",X"4C",X"7E",X"D0",X"01",
		X"34",X"10",X"8E",X"EE",X"65",X"20",X"05",X"34",X"10",X"8E",X"EE",X"73",X"86",X"00",X"BD",X"D0",
		X"55",X"31",X"84",X"35",X"10",X"AF",X"27",X"CC",X"00",X"00",X"ED",X"06",X"ED",X"88",X"10",X"CC",
		X"ED",X"70",X"ED",X"08",X"CC",X"D4",X"DF",X"BD",X"D5",X"4D",X"7E",X"D0",X"0A",X"97",X"73",X"F6",
		X"A1",X"06",X"03",X"AA",X"2B",X"01",X"50",X"D7",X"74",X"8E",X"F2",X"F7",X"86",X"00",X"BD",X"D0",
		X"3E",X"33",X"84",X"96",X"73",X"A7",X"4F",X"4F",X"5F",X"ED",X"47",X"ED",X"49",X"ED",X"4B",X"ED",
		X"4D",X"BD",X"D0",X"95",X"F9",X"29",X"F3",X"BC",X"88",X"88",X"D6",X"74",X"1D",X"ED",X"0E",X"4F",
		X"5F",X"ED",X"88",X"10",X"96",X"73",X"44",X"56",X"9B",X"73",X"D3",X"CC",X"8B",X"80",X"ED",X"0A",
		X"86",X"50",X"A7",X"0C",X"A7",X"C8",X"10",X"EF",X"06",X"9F",X"65",X"96",X"73",X"48",X"8B",X"05",
		X"AF",X"C6",X"0A",X"73",X"26",X"CB",X"39",X"96",X"DF",X"84",X"06",X"8B",X"07",X"AE",X"C6",X"10",
		X"27",X"00",X"B1",X"D6",X"DF",X"86",X"0A",X"C4",X"3F",X"CB",X"E0",X"2B",X"01",X"40",X"10",X"AE",
		X"02",X"31",X"A6",X"10",X"8C",X"F9",X"29",X"24",X"04",X"10",X"8E",X"F9",X"29",X"10",X"8C",X"F9",
		X"47",X"23",X"04",X"10",X"8E",X"F9",X"47",X"10",X"AF",X"02",X"1D",X"E3",X"88",X"10",X"ED",X"88",
		X"10",X"58",X"49",X"58",X"49",X"58",X"49",X"1F",X"89",X"50",X"1D",X"E3",X"88",X"10",X"ED",X"88",
		X"10",X"A6",X"05",X"26",X"3B",X"96",X"DF",X"81",X"40",X"22",X"16",X"84",X"03",X"8B",X"FE",X"AB",
		X"C8",X"10",X"81",X"40",X"24",X"02",X"86",X"40",X"81",X"68",X"25",X"02",X"86",X"68",X"A7",X"C8",
		X"10",X"A6",X"C8",X"10",X"A0",X"0C",X"8B",X"10",X"81",X"20",X"23",X"48",X"80",X"10",X"2B",X"05",
		X"CC",X"FF",X"F0",X"20",X"03",X"CC",X"00",X"10",X"E3",X"88",X"10",X"ED",X"88",X"10",X"20",X"34",
		X"90",X"C0",X"2B",X"12",X"81",X"20",X"25",X"05",X"CC",X"FF",X"F0",X"20",X"19",X"81",X"10",X"22",
		X"1B",X"CC",X"00",X"10",X"20",X"10",X"81",X"E0",X"2E",X"05",X"CC",X"00",X"10",X"20",X"07",X"81",
		X"F0",X"2D",X"09",X"CC",X"FF",X"F0",X"E3",X"88",X"10",X"ED",X"88",X"10",X"96",X"E1",X"84",X"07",
		X"26",X"02",X"8D",X"28",X"86",X"01",X"8E",X"F2",X"F7",X"7E",X"D0",X"01",X"BD",X"F4",X"1D",X"01",
		X"25",X"D5",X"02",X"7A",X"A1",X"13",X"EE",X"06",X"31",X"47",X"AC",X"A1",X"26",X"FC",X"4F",X"5F",
		X"ED",X"3E",X"6A",X"4F",X"26",X"05",X"30",X"C4",X"BD",X"D0",X"15",X"39",X"96",X"99",X"81",X"0A",
		X"24",X"18",X"BD",X"E3",X"F3",X"E4",X"98",X"F9",X"5B",X"E5",X"1E",X"27",X"0D",X"D6",X"E0",X"1D",
		X"58",X"49",X"96",X"DF",X"84",X"1F",X"4C",X"A7",X"88",X"15",X"39",X"BD",X"D0",X"C7",X"34",X"76",
		X"BD",X"F5",X"03",X"EC",X"04",X"10",X"AE",X"02",X"AD",X"B8",X"08",X"35",X"F6",X"34",X"10",X"BD",
		X"D0",X"13",X"35",X"10",X"20",X"0A",X"34",X"10",X"BD",X"D0",X"13",X"35",X"10",X"BD",X"D0",X"C7",
		X"34",X"46",X"EE",X"64",X"37",X"06",X"BD",X"D3",X"60",X"8D",X"09",X"37",X"06",X"EF",X"64",X"BD",
		X"D5",X"4D",X"35",X"C6",X"34",X"76",X"8D",X"C6",X"BD",X"FC",X"63",X"35",X"F6",X"8E",X"F4",X"5B",
		X"AF",X"47",X"86",X"06",X"8E",X"F4",X"4A",X"7E",X"D0",X"01",X"AE",X"47",X"EC",X"81",X"DD",X"33",
		X"A6",X"80",X"97",X"35",X"8C",X"F4",X"64",X"25",X"E7",X"20",X"E2",X"81",X"81",X"2F",X"81",X"2F",
		X"07",X"2F",X"81",X"07",X"86",X"FF",X"97",X"30",X"0F",X"32",X"86",X"03",X"8E",X"F4",X"72",X"7E",
		X"D0",X"01",X"96",X"DF",X"84",X"1F",X"8E",X"E7",X"99",X"A6",X"86",X"97",X"30",X"97",X"32",X"8E",
		X"CC",X"B0",X"9C",X"A6",X"26",X"03",X"8E",X"CC",X"BC",X"9F",X"A6",X"86",X"06",X"8E",X"F4",X"64",
		X"7E",X"D0",X"01",X"96",X"8A",X"26",X"24",X"8E",X"0F",X"1C",X"96",X"8B",X"4A",X"27",X"03",X"8E",
		X"71",X"1C",X"CC",X"18",X"08",X"BD",X"F5",X"C7",X"86",X"08",X"8E",X"F4",X"B0",X"7E",X"D0",X"01",
		X"BD",X"D3",X"D9",X"86",X"0C",X"8E",X"F4",X"93",X"7E",X"D0",X"01",X"7E",X"D0",X"0A",X"DE",X"63",
		X"AF",X"4D",X"D6",X"36",X"E7",X"4C",X"8E",X"F4",X"CC",X"7E",X"D0",X"01",X"A6",X"4C",X"8D",X"3D",
		X"6E",X"D8",X"0D",X"32",X"7D",X"34",X"42",X"96",X"36",X"A7",X"65",X"EE",X"66",X"A6",X"42",X"EE",
		X"C4",X"EF",X"63",X"8D",X"28",X"35",X"42",X"AD",X"F4",X"34",X"42",X"A6",X"65",X"8D",X"1E",X"EE",
		X"66",X"33",X"43",X"EF",X"66",X"35",X"42",X"32",X"63",X"39",X"8D",X"03",X"7E",X"C0",X"00",X"86",
		X"07",X"20",X"0A",X"86",X"02",X"20",X"06",X"86",X"03",X"20",X"02",X"86",X"01",X"97",X"36",X"B7",
		X"D0",X"00",X"39",X"34",X"7F",X"8D",X"EC",X"BD",X"C0",X"02",X"35",X"FF",X"8D",X"E9",X"7E",X"C0",
		X"0F",X"39",X"34",X"76",X"1F",X"01",X"96",X"36",X"34",X"02",X"86",X"02",X"97",X"36",X"B7",X"D0",
		X"00",X"EC",X"A4",X"10",X"AE",X"22",X"34",X"06",X"C5",X"01",X"26",X"17",X"C0",X"02",X"EE",X"A5",
		X"EF",X"85",X"C0",X"02",X"2A",X"F8",X"E6",X"61",X"30",X"89",X"01",X"00",X"31",X"A5",X"4A",X"26",
		X"EB",X"20",X"1D",X"5A",X"A6",X"A5",X"A7",X"85",X"C0",X"02",X"2B",X"08",X"EE",X"A5",X"EF",X"85",
		X"C0",X"02",X"2A",X"F8",X"E6",X"61",X"30",X"89",X"01",X"00",X"31",X"A5",X"6A",X"E4",X"26",X"E3",
		X"32",X"62",X"35",X"02",X"97",X"36",X"B7",X"D0",X"00",X"35",X"F6",X"34",X"56",X"1F",X"01",X"96",
		X"36",X"34",X"02",X"86",X"02",X"97",X"36",X"B7",X"D0",X"00",X"EC",X"A4",X"CE",X"00",X"00",X"34",
		X"04",X"C5",X"01",X"26",X"13",X"C0",X"02",X"EF",X"85",X"C0",X"02",X"2A",X"FA",X"E6",X"E4",X"30",
		X"89",X"01",X"00",X"4A",X"26",X"EF",X"20",X"16",X"5A",X"6F",X"85",X"C0",X"02",X"2B",X"06",X"EF",
		X"85",X"C0",X"02",X"2A",X"FA",X"E6",X"E4",X"30",X"89",X"01",X"00",X"4A",X"26",X"EA",X"35",X"06",
		X"D7",X"36",X"F7",X"D0",X"00",X"35",X"D6",X"34",X"56",X"96",X"36",X"34",X"02",X"A6",X"61",X"20",
		X"BB",X"34",X"76",X"CE",X"9C",X"00",X"8E",X"00",X"00",X"1F",X"12",X"1F",X"10",X"36",X"36",X"36",
		X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"36",X"10",X"11",X"83",X"00",X"00",X"26",X"EE",X"35",
		X"F6",X"34",X"7E",X"CE",X"9C",X"00",X"8E",X"00",X"00",X"1F",X"12",X"1F",X"10",X"1F",X"8B",X"C6",
		X"08",X"36",X"3A",X"36",X"3A",X"36",X"3A",X"36",X"3A",X"5A",X"26",X"F5",X"36",X"3A",X"36",X"3A",
		X"36",X"3A",X"36",X"30",X"33",X"C8",X"D6",X"11",X"83",X"00",X"00",X"26",X"E2",X"35",X"FE",X"7F",
		X"D0",X"00",X"8E",X"CC",X"00",X"6F",X"01",X"6F",X"03",X"6F",X"05",X"6F",X"07",X"86",X"C0",X"A7",
		X"84",X"86",X"FF",X"A7",X"02",X"6F",X"04",X"6F",X"06",X"86",X"04",X"A7",X"03",X"A7",X"05",X"A7",
		X"07",X"8A",X"10",X"A7",X"01",X"8E",X"C0",X"00",X"86",X"C0",X"A7",X"80",X"C6",X"B5",X"3D",X"8C",
		X"C0",X"10",X"26",X"F6",X"1A",X"80",X"1C",X"EF",X"10",X"8E",X"00",X"02",X"4F",X"1F",X"8B",X"1C",
		X"BF",X"5F",X"1F",X"03",X"8E",X"00",X"00",X"53",X"C5",X"09",X"26",X"05",X"53",X"46",X"56",X"20",
		X"0B",X"53",X"C5",X"09",X"26",X"04",X"46",X"56",X"20",X"02",X"44",X"56",X"ED",X"81",X"1E",X"10",
		X"5D",X"26",X"17",X"C6",X"38",X"F7",X"C3",X"FC",X"1F",X"A9",X"C5",X"10",X"27",X"0B",X"7F",X"D0",
		X"00",X"F6",X"CC",X"00",X"53",X"C5",X"03",X"27",X"51",X"5F",X"1E",X"10",X"8C",X"C0",X"00",X"26",
		X"C6",X"1F",X"30",X"8E",X"00",X"00",X"53",X"C5",X"09",X"26",X"05",X"53",X"46",X"56",X"20",X"0B",
		X"53",X"C5",X"09",X"26",X"04",X"46",X"56",X"20",X"02",X"44",X"56",X"10",X"A3",X"81",X"27",X"17",
		X"1E",X"02",X"1F",X"A8",X"85",X"10",X"27",X"0A",X"86",X"03",X"97",X"36",X"B7",X"D0",X"00",X"7E",
		X"C0",X"2A",X"4F",X"1E",X"20",X"1A",X"40",X"1E",X"10",X"5D",X"26",X"42",X"1F",X"A9",X"C5",X"10",
		X"27",X"12",X"F6",X"CC",X"00",X"53",X"C5",X"03",X"26",X"2E",X"86",X"03",X"97",X"36",X"B7",X"D0",
		X"00",X"7E",X"C0",X"2D",X"1F",X"A9",X"C5",X"40",X"27",X"1E",X"1C",X"BF",X"1F",X"B9",X"1F",X"8B",
		X"80",X"03",X"24",X"FC",X"4C",X"26",X"04",X"CA",X"02",X"20",X"09",X"4C",X"26",X"04",X"CA",X"01",
		X"20",X"02",X"CA",X"04",X"1F",X"B8",X"1F",X"9B",X"C6",X"38",X"F7",X"C3",X"FC",X"5F",X"1E",X"10",
		X"8C",X"C0",X"00",X"10",X"26",X"FF",X"7F",X"31",X"3F",X"10",X"26",X"FF",X"35",X"1F",X"A9",X"5D",
		X"2B",X"0B",X"C6",X"03",X"F7",X"D0",X"00",X"BD",X"F8",X"00",X"7E",X"C0",X"30",X"C5",X"10",X"10",
		X"26",X"FF",X"1F",X"86",X"9E",X"1F",X"B9",X"5D",X"27",X"04",X"4C",X"54",X"25",X"FC",X"1F",X"8B",
		X"8B",X"01",X"5F",X"1F",X"04",X"BD",X"F8",X"00",X"CE",X"F8",X"6E",X"7F",X"D0",X"00",X"86",X"38",
		X"B7",X"C3",X"FC",X"A6",X"C4",X"E6",X"C4",X"27",X"2A",X"C4",X"0F",X"F7",X"D0",X"00",X"84",X"70",
		X"44",X"8B",X"C0",X"5F",X"1F",X"01",X"10",X"8E",X"08",X"00",X"1F",X"30",X"C0",X"6C",X"54",X"4F",
		X"E9",X"80",X"31",X"3F",X"26",X"FA",X"C1",X"80",X"27",X"09",X"1F",X"A8",X"85",X"10",X"27",X"3E",
		X"7E",X"F5",X"07",X"33",X"41",X"11",X"83",X"F8",X"86",X"26",X"C0",X"1F",X"A8",X"85",X"10",X"26",
		X"EF",X"1F",X"B8",X"81",X"9E",X"26",X"08",X"BD",X"F5",X"07",X"BD",X"C0",X"00",X"20",X"26",X"C6",
		X"40",X"8D",X"05",X"BD",X"C0",X"03",X"20",X"1D",X"8E",X"CC",X"00",X"E7",X"84",X"E7",X"02",X"7F",
		X"D0",X"00",X"86",X"38",X"B7",X"C3",X"FC",X"30",X"1F",X"26",X"F7",X"7E",X"F5",X"07",X"C6",X"80",
		X"8D",X"E6",X"BD",X"C0",X"06",X"BD",X"C0",X"09",X"7E",X"D7",X"38",X"34",X"03",X"96",X"36",X"34",
		X"02",X"0F",X"36",X"7F",X"D0",X"00",X"E7",X"84",X"35",X"02",X"97",X"36",X"B7",X"D0",X"00",X"35",
		X"83",X"34",X"03",X"96",X"36",X"34",X"02",X"0F",X"36",X"7F",X"D0",X"00",X"E6",X"84",X"20",X"E8",
		X"34",X"06",X"0F",X"52",X"0F",X"49",X"86",X"03",X"97",X"36",X"97",X"48",X"CC",X"FF",X"FF",X"DD",
		X"59",X"35",X"86",X"A6",X"01",X"84",X"0F",X"34",X"02",X"A6",X"81",X"48",X"48",X"48",X"48",X"AB",
		X"E0",X"39",X"34",X"04",X"D6",X"36",X"34",X"04",X"0F",X"36",X"7F",X"D0",X"00",X"8D",X"E4",X"35",
		X"04",X"D7",X"36",X"F7",X"D0",X"00",X"35",X"84",X"8D",X"E8",X"34",X"02",X"8D",X"E4",X"1F",X"89",
		X"35",X"82",X"34",X"02",X"A7",X"01",X"44",X"44",X"44",X"44",X"A7",X"81",X"35",X"82",X"34",X"04",
		X"D6",X"36",X"34",X"04",X"0F",X"36",X"7F",X"D0",X"00",X"8D",X"E7",X"35",X"04",X"D7",X"36",X"F7",
		X"D0",X"00",X"35",X"84",X"8D",X"E8",X"34",X"02",X"1F",X"98",X"8D",X"E2",X"35",X"82",X"20",X"00",
		X"40",X"50",X"60",X"70",X"30",X"00",X"00",X"00",X"07",X"00",X"03",X"00",X"02",X"00",X"01",X"00",
		X"13",X"00",X"12",X"00",X"11",X"00",X"E5",X"91",X"00",X"E8",X"00",X"00",X"00",X"00",X"E8",X"C1",
		X"00",X"F8",X"E9",X"1F",X"00",X"F8",X"D8",X"4E",X"00",X"00",X"D8",X"39",X"00",X"00",X"E8",X"97",
		X"00",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"4C",X"00",X"00",X"D4",X"75",
		X"02",X"00",X"D4",X"3D",X"00",X"00",X"D4",X"6E",X"02",X"00",X"D4",X"7C",X"02",X"00",X"00",X"00",
		X"07",X"28",X"2F",X"81",X"A4",X"15",X"C7",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"08",
		X"F9",X"FB",X"FA",X"23",X"D1",X"93",X"D1",X"1F",X"04",X"08",X"FA",X"4B",X"FA",X"4B",X"D1",X"39",
		X"D1",X"6B",X"04",X"08",X"FA",X"6B",X"FA",X"6B",X"D1",X"39",X"D1",X"6B",X"01",X"01",X"F8",X"F6",
		X"F8",X"F6",X"D8",X"DB",X"D8",X"DB",X"00",X"04",X"08",X"FA",X"8B",X"FA",X"AB",X"D1",X"39",X"D1",
		X"6B",X"02",X"08",X"FA",X"CB",X"FA",X"DB",X"D0",X"F9",X"D1",X"0B",X"02",X"08",X"FA",X"EB",X"FA",
		X"FB",X"D0",X"F9",X"D1",X"0B",X"02",X"08",X"FB",X"0B",X"FB",X"1B",X"D0",X"F9",X"D1",X"0B",X"02",
		X"08",X"FB",X"2B",X"FB",X"3B",X"D0",X"F9",X"D1",X"0B",X"04",X"08",X"FB",X"4B",X"FB",X"6B",X"D1",
		X"39",X"D1",X"6B",X"04",X"08",X"FB",X"8B",X"FB",X"AB",X"D1",X"39",X"D1",X"6B",X"04",X"08",X"FB",
		X"CB",X"FB",X"EB",X"D1",X"39",X"D1",X"6B",X"04",X"08",X"FC",X"0B",X"FC",X"2B",X"D1",X"39",X"D1",
		X"6B",X"04",X"08",X"CC",X"90",X"CC",X"90",X"D1",X"39",X"D1",X"6B",X"02",X"03",X"CC",X"B0",X"CC",
		X"B6",X"D1",X"F1",X"D2",X"0D",X"02",X"03",X"CC",X"BC",X"CC",X"C2",X"D1",X"F1",X"D2",X"0D",X"08",
		X"01",X"F9",X"73",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"03",X"04",X"CC",X"C8",X"CC",
		X"D4",X"D1",X"AD",X"D1",X"D7",X"05",X"08",X"CC",X"E0",X"CD",X"08",X"D1",X"93",X"D1",X"1F",X"05",
		X"08",X"CD",X"30",X"CD",X"58",X"D1",X"93",X"D1",X"1F",X"05",X"08",X"CD",X"80",X"CD",X"A8",X"D1",
		X"93",X"D1",X"1F",X"06",X"04",X"CD",X"D0",X"CD",X"E8",X"D2",X"1F",X"D2",X"60",X"06",X"04",X"CE",
		X"00",X"CE",X"18",X"D2",X"1F",X"D2",X"60",X"06",X"04",X"CE",X"30",X"CE",X"48",X"D2",X"1F",X"D2",
		X"60",X"08",X"06",X"CE",X"60",X"CE",X"90",X"D2",X"8E",X"D2",X"DF",X"08",X"06",X"CE",X"C0",X"CE",
		X"F0",X"D2",X"8E",X"D2",X"DF",X"05",X"04",X"CF",X"20",X"03",X"03",X"CF",X"34",X"06",X"06",X"CF",
		X"3D",X"CF",X"61",X"D3",X"3D",X"D3",X"50",X"06",X"06",X"CF",X"85",X"CF",X"A9",X"D3",X"3D",X"D3",
		X"50",X"08",X"06",X"CF",X"CD",X"CF",X"CD",X"F5",X"22",X"F5",X"7B",X"00",X"00",X"03",X"03",X"00",
		X"00",X"03",X"30",X"0C",X"3C",X"0C",X"08",X"38",X"30",X"00",X"00",X"C0",X"C0",X"C8",X"78",X"78",
		X"70",X"70",X"70",X"00",X"30",X"03",X"03",X"30",X"30",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"03",X"30",X"30",X"03",
		X"03",X"30",X"00",X"CC",X"CC",X"CC",X"87",X"87",X"07",X"07",X"07",X"00",X"03",X"80",X"80",X"83",
		X"03",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"30",X"03",X"00",X"00",X"0D",X"6C",X"6C",
		X"0D",X"00",X"00",X"06",X"E6",X"C8",X"83",X"82",X"C8",X"EC",X"06",X"60",X"6D",X"8C",X"28",X"28",
		X"8C",X"6D",X"60",X"00",X"00",X"E0",X"C6",X"C6",X"E0",X"00",X"00",X"00",X"00",X"02",X"22",X"24",
		X"02",X"00",X"00",X"02",X"22",X"44",X"44",X"24",X"42",X"22",X"00",X"20",X"22",X"44",X"44",X"24",
		X"42",X"22",X"00",X"00",X"00",X"20",X"22",X"22",X"20",X"00",X"00",X"00",X"0E",X"00",X"D8",X"00",
		X"0E",X"00",X"00",X"0F",X"08",X"8C",X"C8",X"8C",X"08",X"0F",X"00",X"00",X"0E",X"80",X"C8",X"80",
		X"0E",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"08",X"8C",X"08",X"E0",X"00",X"00",X"F0",X"80",X"C8",X"8C",X"C8",
		X"80",X"F0",X"00",X"00",X"E0",X"00",X"8D",X"00",X"E0",X"00",X"00",X"33",X"43",X"43",X"87",X"87",
		X"07",X"07",X"07",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"03",X"04",X"04",X"08",X"08",
		X"00",X"00",X"00",X"30",X"30",X"38",X"78",X"78",X"70",X"70",X"70",X"33",X"43",X"43",X"87",X"87",
		X"77",X"77",X"77",X"00",X"00",X"80",X"80",X"80",X"00",X"00",X"00",X"03",X"04",X"04",X"08",X"08",
		X"07",X"07",X"07",X"30",X"30",X"38",X"78",X"78",X"70",X"70",X"70",X"03",X"03",X"83",X"87",X"87",
		X"07",X"07",X"07",X"30",X"40",X"40",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"08",
		X"00",X"00",X"00",X"33",X"34",X"34",X"78",X"78",X"70",X"70",X"70",X"03",X"03",X"83",X"87",X"87",
		X"07",X"07",X"07",X"30",X"40",X"40",X"80",X"80",X"70",X"70",X"70",X"00",X"00",X"08",X"08",X"08",
		X"00",X"00",X"00",X"33",X"34",X"34",X"78",X"78",X"77",X"77",X"77",X"08",X"08",X"DD",X"DE",X"DE",
		X"DE",X"DD",X"00",X"88",X"88",X"DD",X"EE",X"FE",X"EE",X"DD",X"00",X"88",X"88",X"D8",X"D8",X"D8",
		X"D0",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0D",X"0D",
		X"0D",X"0D",X"00",X"88",X"88",X"DD",X"EE",X"EF",X"EE",X"DD",X"00",X"88",X"88",X"DD",X"ED",X"ED",
		X"ED",X"DD",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"08",X"DD",X"DE",X"DE",
		X"DE",X"DD",X"00",X"00",X"88",X"DD",X"EE",X"FE",X"EE",X"DD",X"00",X"00",X"88",X"D8",X"D8",X"D8",
		X"D8",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0D",X"0D",
		X"0D",X"0D",X"00",X"00",X"88",X"DD",X"EE",X"EF",X"EE",X"DD",X"00",X"00",X"88",X"DD",X"ED",X"ED",
		X"ED",X"DD",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"DD",X"DE",X"DE",
		X"DE",X"DD",X"00",X"00",X"00",X"DD",X"EE",X"FE",X"EE",X"DD",X"00",X"00",X"00",X"D8",X"D8",X"D8",
		X"D8",X"D8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0D",X"0D",
		X"0D",X"0D",X"00",X"00",X"00",X"DD",X"EE",X"EF",X"EE",X"DD",X"00",X"00",X"00",X"DD",X"ED",X"ED",
		X"ED",X"DD",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"DD",X"DE",X"DE",
		X"DE",X"DD",X"00",X"00",X"00",X"DD",X"EE",X"FE",X"EE",X"DD",X"88",X"00",X"00",X"D0",X"D8",X"D8",
		X"D8",X"D8",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0D",X"0D",
		X"0D",X"0D",X"00",X"00",X"00",X"DD",X"EE",X"EF",X"EE",X"DD",X"88",X"00",X"00",X"DD",X"ED",X"ED",
		X"ED",X"DD",X"88",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"FC",X"69",X"7E",X"FC",X"CC",X"7E",X"FD",X"2D",X"34",X"66",X"EC",X"02",X"34",X"06",X"FC",
		X"FF",X"9D",X"ED",X"02",X"9F",X"65",X"EC",X"0A",X"93",X"20",X"10",X"83",X"26",X"00",X"22",X"17",
		X"10",X"9E",X"E2",X"27",X"09",X"31",X"A8",X"40",X"10",X"8C",X"A0",X"00",X"26",X"04",X"10",X"8E",
		X"9C",X"00",X"10",X"9C",X"E2",X"26",X"06",X"35",X"06",X"ED",X"02",X"20",X"2D",X"A6",X"A4",X"2B",
		X"E4",X"27",X"03",X"BD",X"FD",X"D5",X"96",X"BA",X"85",X"80",X"26",X"06",X"FC",X"FF",X"DD",X"BD",
		X"FF",X"DA",X"A6",X"88",X"14",X"8A",X"02",X"A7",X"88",X"14",X"CC",X"AF",X"00",X"ED",X"A4",X"35",
		X"06",X"ED",X"22",X"33",X"A8",X"40",X"EF",X"24",X"AF",X"2A",X"35",X"E6",X"34",X"66",X"EC",X"0A",
		X"93",X"20",X"81",X"26",X"22",X"55",X"DD",X"E9",X"10",X"9E",X"E2",X"27",X"09",X"31",X"A8",X"40",
		X"10",X"8C",X"A0",X"00",X"26",X"04",X"10",X"8E",X"9C",X"00",X"10",X"9C",X"E2",X"27",X"3C",X"A6",
		X"A4",X"2B",X"EA",X"27",X"03",X"BD",X"FD",X"D5",X"10",X"9F",X"E2",X"CC",X"01",X"00",X"ED",X"A4",
		X"EC",X"02",X"ED",X"22",X"33",X"A8",X"40",X"EF",X"24",X"DC",X"E9",X"58",X"49",X"58",X"49",X"E6",
		X"0C",X"ED",X"28",X"93",X"F8",X"EE",X"22",X"AB",X"C4",X"24",X"08",X"EB",X"41",X"24",X"04",X"DC",
		X"F8",X"20",X"06",X"EC",X"C4",X"44",X"54",X"E3",X"28",X"ED",X"26",X"35",X"E6",X"10",X"8E",X"9C",
		X"00",X"96",X"BA",X"85",X"04",X"27",X"0C",X"A6",X"A4",X"2B",X"56",X"CC",X"00",X"00",X"ED",X"A4",
		X"7E",X"FD",X"C9",X"EC",X"A4",X"10",X"27",X"00",X"80",X"2B",X"33",X"C3",X"00",X"AA",X"ED",X"A4",
		X"81",X"30",X"23",X"0A",X"BD",X"FD",X"D5",X"CC",X"00",X"00",X"ED",X"A4",X"20",X"6B",X"DC",X"20",
		X"C4",X"C0",X"34",X"06",X"DC",X"22",X"C4",X"C0",X"A3",X"E1",X"58",X"49",X"58",X"49",X"34",X"02",
		X"A6",X"26",X"AB",X"E4",X"A7",X"26",X"A6",X"28",X"AB",X"E0",X"A7",X"28",X"20",X"45",X"83",X"01",
		X"00",X"ED",X"A4",X"2A",X"0C",X"AE",X"2A",X"EC",X"0A",X"93",X"20",X"8B",X"0C",X"85",X"C0",X"27",
		X"18",X"CC",X"00",X"00",X"ED",X"A4",X"EC",X"22",X"AE",X"2A",X"ED",X"02",X"A6",X"88",X"14",X"84",
		X"FD",X"A7",X"88",X"14",X"BD",X"FD",X"D5",X"20",X"20",X"80",X"0C",X"58",X"49",X"58",X"49",X"E6",
		X"0C",X"ED",X"28",X"C6",X"DA",X"3D",X"48",X"EE",X"22",X"E6",X"C4",X"3D",X"E6",X"41",X"54",X"E3",
		X"28",X"ED",X"26",X"BD",X"FD",X"D5",X"BD",X"FD",X"EF",X"31",X"A8",X"40",X"10",X"8C",X"A0",X"00",
		X"10",X"26",X"FF",X"5D",X"39",X"34",X"16",X"CC",X"00",X"00",X"30",X"A8",X"40",X"9F",X"F3",X"AE",
		X"24",X"9C",X"F3",X"27",X"08",X"ED",X"91",X"9C",X"F3",X"26",X"FA",X"AF",X"24",X"35",X"96",X"34",
		X"76",X"10",X"9F",X"F6",X"A6",X"A4",X"84",X"7F",X"97",X"E7",X"33",X"A8",X"40",X"0F",X"E6",X"AE",
		X"22",X"EC",X"02",X"DD",X"F3",X"EC",X"84",X"97",X"F1",X"D7",X"F2",X"C5",X"01",X"26",X"05",X"8E",
		X"FF",X"27",X"20",X"03",X"8E",X"FE",X"F3",X"9F",X"ED",X"EC",X"26",X"A3",X"28",X"97",X"E4",X"54",
		X"D7",X"E5",X"09",X"E6",X"96",X"E7",X"D6",X"E4",X"3D",X"DD",X"E9",X"E6",X"26",X"4F",X"93",X"E9",
		X"DD",X"E9",X"4D",X"27",X"18",X"DC",X"F3",X"DB",X"F2",X"89",X"00",X"DD",X"F3",X"0A",X"F1",X"10",
		X"27",X"00",X"F2",X"DC",X"E9",X"DB",X"E7",X"89",X"00",X"DD",X"E9",X"20",X"E5",X"C1",X"98",X"10",
		X"22",X"00",X"E2",X"96",X"E7",X"48",X"97",X"E8",X"D6",X"E5",X"3D",X"DD",X"EB",X"E6",X"27",X"4F",
		X"93",X"EB",X"D0",X"E6",X"89",X"00",X"0F",X"F5",X"4D",X"26",X"04",X"C1",X"2A",X"24",X"10",X"0C",
		X"F5",X"0A",X"F2",X"0A",X"F2",X"10",X"2F",X"00",X"BC",X"DB",X"E8",X"89",X"00",X"20",X"E9",X"DD",
		X"EB",X"96",X"F2",X"84",X"FE",X"8E",X"FF",X"48",X"AE",X"86",X"9F",X"EF",X"9E",X"F3",X"08",X"F5",
		X"96",X"EA",X"D6",X"F5",X"3A",X"D6",X"EC",X"6E",X"9F",X"A0",X"EF",X"ED",X"C3",X"10",X"AE",X"81",
		X"10",X"AF",X"D4",X"DB",X"E8",X"25",X"56",X"ED",X"C3",X"10",X"AE",X"81",X"10",X"AF",X"D4",X"DB",
		X"E8",X"25",X"50",X"ED",X"C3",X"10",X"AE",X"81",X"10",X"AF",X"D4",X"DB",X"E8",X"25",X"4A",X"ED",
		X"C3",X"10",X"AE",X"81",X"10",X"AF",X"D4",X"DB",X"E8",X"25",X"44",X"ED",X"C3",X"10",X"AE",X"81",
		X"10",X"AF",X"D4",X"DB",X"E8",X"25",X"3E",X"ED",X"C3",X"10",X"AE",X"81",X"10",X"AF",X"D4",X"DB",
		X"E8",X"25",X"38",X"ED",X"C3",X"10",X"AE",X"81",X"10",X"AF",X"D4",X"DB",X"E8",X"25",X"32",X"6E",
		X"9F",X"A0",X"ED",X"25",X"30",X"ED",X"C3",X"E6",X"80",X"E7",X"D4",X"20",X"2A",X"30",X"0C",X"6E",
		X"9F",X"A0",X"ED",X"30",X"0A",X"6E",X"9F",X"A0",X"ED",X"30",X"08",X"6E",X"9F",X"A0",X"ED",X"30",
		X"06",X"6E",X"9F",X"A0",X"ED",X"30",X"04",X"6E",X"9F",X"A0",X"ED",X"30",X"02",X"6E",X"9F",X"A0",
		X"ED",X"6E",X"9F",X"A0",X"ED",X"30",X"01",X"0A",X"F1",X"27",X"0A",X"9B",X"E7",X"25",X"06",X"81",
		X"98",X"10",X"23",X"FF",X"5D",X"9E",X"F6",X"EF",X"04",X"EC",X"06",X"81",X"98",X"22",X"07",X"D0",
		X"E6",X"8E",X"00",X"00",X"AF",X"8B",X"35",X"F6",X"FE",X"EF",X"FE",X"E3",X"FE",X"D7",X"FE",X"CB",
		X"FE",X"BF",X"FE",X"B3",X"FE",X"A7",X"FE",X"9B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"EC",X"F8",
		X"6E",X"7E",X"F8",X"22",X"7E",X"F8",X"3A",X"7E",X"F8",X"38",X"7E",X"F8",X"4E",X"7E",X"F8",X"66",
		X"7E",X"F8",X"64",X"7E",X"F5",X"22",X"7E",X"F5",X"7B",X"7E",X"F5",X"C7",X"7E",X"F5",X"D1",X"7E",
		X"F7",X"58",X"7E",X"F7",X"93",X"7E",X"F6",X"62",X"7E",X"F7",X"D5",X"7E",X"F4",X"FA",X"7E",X"F4",
		X"D3",X"7E",X"F4",X"BE",X"7E",X"F7",X"DB",X"7E",X"F7",X"F1",X"7E",X"D5",X"4D",X"D4",X"EE",X"2A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F6",X"1F",X"F6",X"1F",X"F6",X"1F",X"F6",X"1F",X"A0",X"8F",X"F6",X"1F",X"F6",X"1F",X"F6",X"1F",
		X"7E",X"C0",X"06",X"7E",X"CC",X"AD",X"BD",X"D0",X"7C",X"86",X"FF",X"97",X"BA",X"BD",X"E0",X"52",
		X"96",X"37",X"B7",X"A1",X"83",X"4F",X"B7",X"A1",X"84",X"B7",X"A1",X"78",X"96",X"B7",X"10",X"27",
		X"06",X"55",X"8E",X"C8",X"F4",X"86",X"00",X"BD",X"D0",X"55",X"10",X"8E",X"A1",X"C2",X"86",X"01",
		X"97",X"06",X"10",X"BF",X"A1",X"7B",X"8E",X"B2",X"B4",X"BD",X"C1",X"47",X"10",X"24",X"00",X"EA",
		X"7C",X"A1",X"78",X"BD",X"F5",X"D1",X"96",X"06",X"4A",X"26",X"05",X"BD",X"D8",X"DC",X"20",X"03",
		X"BD",X"D8",X"EA",X"C6",X"85",X"D7",X"27",X"86",X"3E",X"8E",X"B2",X"60",X"BD",X"C1",X"47",X"24",
		X"02",X"86",X"3D",X"8E",X"CC",X"02",X"C6",X"3F",X"BD",X"FF",X"D4",X"C6",X"24",X"BD",X"FF",X"D4",
		X"5A",X"26",X"FD",X"C6",X"3F",X"BD",X"FF",X"D4",X"1F",X"89",X"BD",X"FF",X"D4",X"CE",X"C0",X"ED",
		X"96",X"06",X"48",X"33",X"C6",X"8E",X"3E",X"38",X"BD",X"FF",X"CE",X"C0",X"02",X"02",X"CE",X"C0",
		X"FD",X"8E",X"14",X"58",X"BD",X"FF",X"CE",X"C0",X"02",X"02",X"CC",X"41",X"2F",X"DD",X"00",X"86",
		X"40",X"DD",X"02",X"DD",X"04",X"BD",X"C1",X"58",X"86",X"28",X"B7",X"A1",X"7D",X"8E",X"C1",X"DC",
		X"86",X"00",X"BD",X"D0",X"55",X"8E",X"C1",X"E7",X"86",X"00",X"BD",X"D0",X"55",X"8E",X"C1",X"FA",
		X"86",X"00",X"BD",X"D0",X"55",X"7F",X"A1",X"7A",X"BD",X"C1",X"6B",X"4F",X"B7",X"A1",X"86",X"B7",
		X"A1",X"85",X"86",X"01",X"8E",X"C0",X"DA",X"7E",X"F4",X"BE",X"96",X"7B",X"85",X"01",X"26",X"14",
		X"7D",X"A1",X"7D",X"27",X"29",X"7C",X"A1",X"86",X"B6",X"A1",X"86",X"81",X"05",X"26",X"E3",X"B7",
		X"A1",X"85",X"20",X"DE",X"7F",X"A1",X"86",X"7D",X"A1",X"85",X"27",X"D6",X"86",X"14",X"B7",X"A1",
		X"7D",X"7C",X"A1",X"7A",X"BD",X"C1",X"6B",X"B6",X"A1",X"7A",X"81",X"03",X"26",X"BD",X"BD",X"D0",
		X"7C",X"8E",X"B2",X"A8",X"CE",X"B2",X"54",X"BD",X"C1",X"94",X"8E",X"C4",X"71",X"8D",X"28",X"24",
		X"09",X"8E",X"C4",X"65",X"CE",X"C4",X"11",X"BD",X"C1",X"94",X"10",X"8E",X"A1",X"FF",X"96",X"06",
		X"4C",X"81",X"03",X"10",X"26",X"FE",X"F9",X"7D",X"A1",X"78",X"26",X"08",X"86",X"FF",X"8E",X"C1",
		X"44",X"7E",X"F4",X"BE",X"7E",X"C2",X"63",X"34",X"16",X"BD",X"F8",X"38",X"10",X"A3",X"21",X"26",
		X"05",X"BD",X"F8",X"22",X"A1",X"23",X"35",X"96",X"8E",X"46",X"AC",X"CC",X"14",X"08",X"BD",X"F5",
		X"C7",X"CE",X"C0",X"FF",X"BD",X"FF",X"CE",X"C0",X"02",X"02",X"39",X"7F",X"A1",X"62",X"8E",X"45",
		X"B7",X"CE",X"11",X"11",X"B6",X"A1",X"62",X"B1",X"A1",X"7A",X"26",X"03",X"CE",X"DD",X"DD",X"CC",
		X"04",X"00",X"EF",X"8B",X"4A",X"26",X"FB",X"7C",X"A1",X"62",X"30",X"89",X"08",X"00",X"8C",X"5D",
		X"B7",X"26",X"DE",X"39",X"FF",X"A1",X"64",X"10",X"BE",X"A1",X"7B",X"8D",X"AA",X"24",X"09",X"8D",
		X"24",X"30",X"14",X"BC",X"A1",X"64",X"22",X"F3",X"30",X"0C",X"EC",X"21",X"BD",X"F8",X"64",X"A6",
		X"23",X"BD",X"F8",X"4E",X"CE",X"A0",X"00",X"A6",X"C4",X"BD",X"F8",X"4E",X"33",X"42",X"11",X"83",
		X"A0",X"06",X"26",X"F3",X"39",X"34",X"10",X"BD",X"F8",X"38",X"30",X"08",X"BD",X"F8",X"64",X"30",
		X"88",X"E8",X"AC",X"E4",X"27",X"04",X"30",X"0C",X"20",X"ED",X"35",X"90",X"7A",X"A1",X"7D",X"86",
		X"3C",X"8E",X"C1",X"DC",X"7E",X"F4",X"BE",X"96",X"33",X"26",X"04",X"96",X"27",X"20",X"01",X"4F",
		X"97",X"33",X"86",X"0F",X"8E",X"C1",X"E7",X"7E",X"F4",X"BE",X"7F",X"A1",X"79",X"96",X"7B",X"85",
		X"80",X"27",X"04",X"86",X"FF",X"20",X"0F",X"96",X"7D",X"85",X"01",X"27",X"04",X"86",X"01",X"20",
		X"05",X"7F",X"A1",X"79",X"20",X"34",X"B1",X"A1",X"79",X"26",X"37",X"7A",X"A1",X"7F",X"26",X"2A",
		X"8E",X"A0",X"00",X"F6",X"A1",X"7A",X"58",X"3A",X"A6",X"84",X"BB",X"A1",X"79",X"81",X"3F",X"26",
		X"02",X"86",X"5A",X"81",X"5B",X"26",X"02",X"86",X"40",X"A7",X"84",X"BD",X"C1",X"58",X"B6",X"A1",
		X"7E",X"44",X"8B",X"05",X"B7",X"A1",X"7E",X"B7",X"A1",X"7F",X"86",X"01",X"8E",X"C1",X"FD",X"7E",
		X"F4",X"BE",X"B7",X"A1",X"79",X"86",X"37",X"B7",X"A1",X"7E",X"86",X"03",X"B7",X"A1",X"7F",X"20",
		X"E9",X"DE",X"FF",X"7F",X"A1",X"62",X"BD",X"D0",X"7C",X"BD",X"C8",X"6F",X"BD",X"F5",X"D1",X"BD",
		X"D8",X"DC",X"0F",X"27",X"8E",X"C8",X"F4",X"86",X"00",X"BD",X"D0",X"55",X"BD",X"C9",X"36",X"CE",
		X"C1",X"01",X"8E",X"38",X"54",X"BD",X"FF",X"CE",X"C0",X"02",X"02",X"CE",X"11",X"11",X"8E",X"1E",
		X"7B",X"CC",X"5F",X"00",X"EF",X"8B",X"81",X"41",X"26",X"02",X"86",X"1F",X"4A",X"2A",X"F5",X"86",
		X"2F",X"97",X"07",X"97",X"0B",X"97",X"12",X"CE",X"C1",X"03",X"8E",X"18",X"86",X"BF",X"A1",X"81",
		X"8E",X"B2",X"60",X"BF",X"A1",X"64",X"8D",X"4E",X"8E",X"59",X"86",X"BF",X"A1",X"81",X"8E",X"C4",
		X"1D",X"BF",X"A1",X"64",X"8D",X"40",X"86",X"3F",X"97",X"32",X"10",X"8E",X"B3",X"00",X"CC",X"3C",
		X"18",X"ED",X"A4",X"CC",X"B4",X"12",X"ED",X"22",X"CC",X"30",X"38",X"BD",X"F5",X"22",X"8E",X"E7",
		X"82",X"86",X"00",X"BD",X"D0",X"55",X"86",X"3C",X"B7",X"A1",X"7D",X"7D",X"A1",X"84",X"26",X"14",
		X"7D",X"A1",X"62",X"10",X"26",X"FF",X"6C",X"7A",X"A1",X"7D",X"27",X"08",X"86",X"0A",X"8E",X"C2",
		X"EB",X"7E",X"F4",X"BE",X"20",X"4B",X"86",X"31",X"97",X"06",X"4F",X"10",X"8E",X"A0",X"0C",X"BE",
		X"A1",X"64",X"BD",X"FF",X"D7",X"30",X"01",X"C4",X"0F",X"26",X"07",X"4D",X"26",X"04",X"C6",X"40",
		X"20",X"03",X"4C",X"CB",X"30",X"E7",X"A0",X"10",X"8C",X"A0",X"12",X"26",X"E5",X"BD",X"F8",X"38",
		X"DD",X"08",X"BD",X"F8",X"22",X"97",X"0A",X"BF",X"A1",X"64",X"BE",X"A1",X"81",X"BD",X"FF",X"CE",
		X"C0",X"02",X"02",X"30",X"0A",X"BF",X"A1",X"81",X"0C",X"06",X"96",X"06",X"81",X"39",X"26",X"BA",
		X"39",X"BD",X"D0",X"7C",X"BD",X"C4",X"3C",X"86",X"D9",X"97",X"BA",X"BD",X"C9",X"36",X"8E",X"C8",
		X"F4",X"86",X"00",X"BD",X"D0",X"55",X"BD",X"D6",X"BC",X"8E",X"CC",X"63",X"BF",X"A1",X"96",X"8E",
		X"E7",X"82",X"86",X"00",X"BD",X"D0",X"55",X"8E",X"F4",X"64",X"86",X"00",X"BD",X"D0",X"55",X"8E",
		X"F4",X"3D",X"86",X"00",X"BD",X"D0",X"55",X"8E",X"E9",X"E3",X"86",X"00",X"BD",X"D0",X"55",X"8E",
		X"C6",X"4F",X"86",X"00",X"BD",X"D0",X"55",X"BD",X"D0",X"AD",X"CC",X"00",X"00",X"ED",X"0E",X"ED",
		X"88",X"10",X"CC",X"1E",X"00",X"ED",X"0A",X"CC",X"DB",X"00",X"ED",X"0C",X"CC",X"F9",X"01",X"ED",
		X"02",X"9F",X"65",X"CC",X"66",X"66",X"ED",X"88",X"12",X"BF",X"A1",X"89",X"BD",X"D0",X"AD",X"CC",
		X"00",X"00",X"ED",X"0E",X"ED",X"88",X"10",X"CC",X"08",X"00",X"ED",X"0A",X"CC",X"50",X"00",X"ED",
		X"0C",X"CC",X"F9",X"C1",X"ED",X"02",X"9F",X"65",X"CC",X"00",X"00",X"ED",X"88",X"12",X"BF",X"A1",
		X"8B",X"BD",X"D0",X"AD",X"CC",X"F9",X"85",X"ED",X"02",X"CC",X"1D",X"A0",X"ED",X"0A",X"CC",X"40",
		X"00",X"ED",X"0C",X"CC",X"00",X"A0",X"ED",X"88",X"10",X"CC",X"00",X"00",X"ED",X"0E",X"CC",X"44",
		X"33",X"ED",X"88",X"12",X"BD",X"FC",X"60",X"BF",X"A1",X"8D",X"86",X"E6",X"8E",X"C4",X"12",X"7E",
		X"F4",X"BE",X"CC",X"FF",X"50",X"BE",X"A1",X"8D",X"ED",X"88",X"10",X"BE",X"A1",X"89",X"ED",X"88",
		X"10",X"86",X"A0",X"8E",X"C4",X"29",X"7E",X"F4",X"BE",X"8E",X"C5",X"F5",X"86",X"00",X"BD",X"D0",
		X"55",X"BF",X"A1",X"87",X"86",X"15",X"8E",X"C4",X"75",X"7E",X"F4",X"BE",X"86",X"FF",X"97",X"BA",
		X"BD",X"D8",X"05",X"BD",X"F5",X"D1",X"CC",X"00",X"00",X"DD",X"20",X"DD",X"22",X"BD",X"FF",X"CE",
		X"F4",X"FA",X"00",X"BD",X"D7",X"F5",X"86",X"DB",X"97",X"BA",X"8E",X"10",X"30",X"9F",X"BF",X"39",
		X"BE",X"A1",X"87",X"FE",X"A1",X"94",X"4F",X"A7",X"C4",X"33",X"C9",X"01",X"00",X"11",X"A3",X"07",
		X"23",X"F5",X"7E",X"D0",X"15",X"8D",X"E9",X"BE",X"A1",X"8D",X"BD",X"D0",X"C7",X"BD",X"FC",X"63",
		X"BE",X"A1",X"8B",X"CC",X"00",X"40",X"ED",X"0E",X"CC",X"00",X"D4",X"ED",X"88",X"10",X"86",X"2D",
		X"B7",X"A1",X"8F",X"BE",X"A1",X"89",X"CC",X"00",X"00",X"ED",X"88",X"10",X"BE",X"A1",X"89",X"EC",
		X"88",X"10",X"C3",X"00",X"08",X"ED",X"88",X"10",X"7A",X"A1",X"8F",X"27",X"08",X"86",X"02",X"8E",
		X"C4",X"9C",X"7E",X"F4",X"BE",X"BD",X"D0",X"AD",X"CC",X"00",X"00",X"ED",X"0E",X"ED",X"88",X"10",
		X"CC",X"1D",X"FF",X"ED",X"0A",X"CC",X"90",X"00",X"ED",X"0C",X"CC",X"F9",X"E7",X"ED",X"02",X"9F",
		X"65",X"CC",X"00",X"00",X"ED",X"88",X"12",X"BF",X"A1",X"90",X"CC",X"00",X"00",X"CE",X"00",X"C0",
		X"BE",X"A1",X"8B",X"ED",X"0E",X"EF",X"88",X"10",X"BE",X"A1",X"89",X"CC",X"1E",X"80",X"ED",X"0A",
		X"CC",X"A2",X"E0",X"ED",X"0C",X"EF",X"88",X"10",X"86",X"50",X"8E",X"C5",X"00",X"7E",X"F4",X"BE",
		X"BE",X"A1",X"90",X"CC",X"E0",X"00",X"ED",X"0C",X"CC",X"1C",X"00",X"ED",X"0A",X"BE",X"A1",X"89",
		X"CC",X"00",X"00",X"ED",X"88",X"10",X"BE",X"A1",X"8B",X"CC",X"F9",X"CB",X"ED",X"02",X"CC",X"FF",
		X"C0",X"ED",X"0E",X"CC",X"FE",X"80",X"ED",X"88",X"10",X"86",X"60",X"8E",X"C5",X"31",X"7E",X"F4",
		X"BE",X"BE",X"A1",X"8B",X"CC",X"F9",X"C1",X"ED",X"02",X"CC",X"00",X"00",X"ED",X"0E",X"ED",X"88",
		X"10",X"BE",X"A1",X"90",X"EC",X"04",X"BD",X"D0",X"C7",X"BD",X"D3",X"50",X"CE",X"CC",X"7D",X"BD",
		X"D0",X"AD",X"EC",X"C9",X"00",X"0C",X"ED",X"02",X"EC",X"C9",X"00",X"24",X"ED",X"88",X"12",X"CC",
		X"1F",X"00",X"ED",X"0A",X"CC",X"A0",X"00",X"ED",X"0C",X"CC",X"FF",X"40",X"ED",X"88",X"10",X"CC",
		X"00",X"00",X"ED",X"0E",X"BD",X"FC",X"60",X"FF",X"A1",X"92",X"BF",X"A1",X"8D",X"86",X"5F",X"8E",
		X"C5",X"85",X"7E",X"F4",X"BE",X"8E",X"C5",X"F5",X"86",X"00",X"BD",X"D0",X"55",X"BF",X"A1",X"87",
		X"86",X"17",X"8E",X"C5",X"98",X"7E",X"F4",X"BE",X"BD",X"C4",X"60",X"BE",X"A1",X"8D",X"BD",X"D0",
		X"C7",X"BD",X"D0",X"AD",X"BD",X"FC",X"63",X"FE",X"A1",X"92",X"EC",X"C9",X"00",X"18",X"ED",X"0A",
		X"EC",X"C1",X"ED",X"0C",X"CC",X"00",X"00",X"ED",X"88",X"10",X"ED",X"0E",X"BD",X"FC",X"60",X"FF",
		X"A1",X"92",X"86",X"20",X"8E",X"C5",X"CA",X"7E",X"F4",X"BE",X"BE",X"A1",X"96",X"30",X"02",X"BF",
		X"A1",X"96",X"86",X"20",X"8E",X"C5",X"DA",X"7E",X"F4",X"BE",X"FE",X"A1",X"92",X"11",X"83",X"CC",
		X"89",X"10",X"26",X"FF",X"6A",X"86",X"FF",X"8E",X"C5",X"ED",X"7E",X"F4",X"BE",X"86",X"FF",X"8E",
		X"C6",X"77",X"7E",X"F4",X"BE",X"BE",X"A1",X"8B",X"AE",X"04",X"30",X"89",X"07",X"04",X"AF",X"47",
		X"AF",X"49",X"BF",X"A1",X"94",X"86",X"04",X"AE",X"47",X"C6",X"11",X"E7",X"84",X"30",X"89",X"01",
		X"00",X"4A",X"26",X"F7",X"C6",X"99",X"E7",X"84",X"AF",X"47",X"10",X"9E",X"A4",X"10",X"8C",X"A1",
		X"5F",X"25",X"04",X"10",X"8E",X"A1",X"42",X"AE",X"49",X"86",X"03",X"E6",X"A0",X"E7",X"84",X"30",
		X"89",X"01",X"00",X"4A",X"26",X"F5",X"10",X"9F",X"A4",X"AF",X"49",X"BE",X"A1",X"94",X"6F",X"84",
		X"30",X"89",X"01",X"00",X"BF",X"A1",X"94",X"86",X"01",X"8E",X"C6",X"05",X"7E",X"F4",X"BE",X"10",
		X"8E",X"CC",X"61",X"EE",X"A9",X"00",X"0E",X"AE",X"A1",X"BD",X"FF",X"CE",X"C0",X"02",X"02",X"10",
		X"BF",X"A1",X"98",X"86",X"06",X"8E",X"C6",X"6B",X"7E",X"F4",X"BE",X"10",X"BE",X"A1",X"98",X"10",
		X"BC",X"A1",X"96",X"26",X"DE",X"20",X"D8",X"BD",X"D0",X"7C",X"7F",X"A1",X"84",X"86",X"FB",X"97",
		X"BA",X"BD",X"F5",X"D1",X"0F",X"52",X"CC",X"FF",X"FF",X"DD",X"59",X"8E",X"E7",X"82",X"86",X"00",
		X"BD",X"D0",X"55",X"8E",X"F4",X"3D",X"86",X"00",X"BD",X"D0",X"55",X"86",X"3F",X"97",X"32",X"7E",
		X"C6",X"A2",X"BD",X"C8",X"6F",X"86",X"03",X"B7",X"A1",X"6A",X"8E",X"C9",X"41",X"BF",X"A1",X"6B",
		X"B6",X"A1",X"6A",X"B7",X"A1",X"63",X"10",X"BE",X"A1",X"6B",X"A6",X"A0",X"81",X"AA",X"23",X"0E",
		X"43",X"27",X"F7",X"4A",X"26",X"4B",X"EC",X"A1",X"FD",X"A1",X"66",X"4F",X"20",X"18",X"48",X"24",
		X"03",X"7A",X"A1",X"66",X"48",X"24",X"03",X"7C",X"A1",X"66",X"48",X"24",X"03",X"7A",X"A1",X"67",
		X"48",X"24",X"03",X"7C",X"A1",X"67",X"B7",X"A1",X"62",X"FC",X"A1",X"66",X"44",X"1F",X"01",X"E6",
		X"84",X"25",X"04",X"CA",X"F0",X"20",X"02",X"CA",X"0F",X"E7",X"84",X"B6",X"A1",X"62",X"26",X"CE",
		X"7A",X"A1",X"63",X"26",X"B5",X"10",X"BF",X"A1",X"6B",X"86",X"02",X"8E",X"C6",X"B0",X"BD",X"F4",
		X"BE",X"BF",X"A1",X"68",X"86",X"03",X"B1",X"A1",X"6A",X"26",X"0D",X"86",X"0A",X"B7",X"A1",X"6A",
		X"8E",X"C7",X"30",X"86",X"00",X"BD",X"D0",X"55",X"8E",X"C9",X"41",X"BF",X"A1",X"6B",X"20",X"80",
		X"8E",X"C7",X"4C",X"86",X"00",X"BD",X"D0",X"55",X"8E",X"32",X"58",X"CE",X"C0",X"ED",X"BD",X"FF",
		X"CE",X"C0",X"02",X"02",X"86",X"05",X"8E",X"C7",X"38",X"BD",X"F4",X"BE",X"86",X"30",X"8E",X"C7",
		X"54",X"7E",X"F4",X"BE",X"CC",X"B3",X"D6",X"FD",X"A1",X"6D",X"CC",X"B4",X"12",X"FD",X"A1",X"6F",
		X"CC",X"00",X"00",X"DD",X"20",X"CC",X"0C",X"00",X"FD",X"A1",X"71",X"CC",X"B3",X"04",X"FD",X"A1",
		X"73",X"BE",X"A1",X"73",X"10",X"BE",X"A1",X"6D",X"CC",X"04",X"0C",X"ED",X"A4",X"FC",X"A1",X"6F",
		X"ED",X"22",X"C3",X"00",X"60",X"FD",X"A1",X"6F",X"10",X"AF",X"02",X"FC",X"A1",X"71",X"ED",X"0A",
		X"C3",X"01",X"00",X"FD",X"A1",X"71",X"CC",X"98",X"00",X"ED",X"0C",X"BD",X"FC",X"60",X"30",X"0E",
		X"BF",X"A1",X"73",X"31",X"24",X"10",X"BF",X"A1",X"6D",X"10",X"8C",X"B4",X"12",X"26",X"C2",X"86",
		X"2E",X"8E",X"C7",X"B7",X"7E",X"F4",X"BE",X"8E",X"B3",X"00",X"CC",X"3C",X"18",X"ED",X"84",X"CC",
		X"B4",X"12",X"ED",X"02",X"8E",X"C8",X"48",X"86",X"00",X"BD",X"D0",X"55",X"86",X"28",X"8E",X"C7",
		X"D4",X"7E",X"F4",X"BE",X"8E",X"F4",X"64",X"86",X"00",X"BD",X"D0",X"55",X"FE",X"A1",X"68",X"10",
		X"8E",X"CC",X"11",X"8E",X"3B",X"D0",X"EC",X"A1",X"FD",X"A1",X"64",X"86",X"01",X"5F",X"B5",X"A1",
		X"64",X"27",X"02",X"C6",X"10",X"B5",X"A1",X"65",X"27",X"02",X"CA",X"01",X"E7",X"80",X"48",X"26",
		X"EC",X"30",X"89",X"00",X"F8",X"10",X"8C",X"CC",X"61",X"26",X"DB",X"8E",X"A0",X"26",X"F6",X"C6",
		X"F8",X"A6",X"85",X"43",X"84",X"07",X"26",X"08",X"8E",X"80",X"18",X"CC",X"20",X"A0",X"EF",X"8B",
		X"86",X"01",X"97",X"B7",X"8E",X"C8",X"F4",X"86",X"00",X"BD",X"D0",X"55",X"86",X"3C",X"B7",X"A1",
		X"7D",X"7D",X"A1",X"84",X"10",X"26",X"FB",X"19",X"7A",X"A1",X"7D",X"27",X"08",X"86",X"0A",X"8E",
		X"C8",X"31",X"7E",X"F4",X"BE",X"7E",X"C2",X"63",X"10",X"8E",X"B3",X"00",X"CC",X"30",X"90",X"BD",
		X"F5",X"22",X"7D",X"9C",X"00",X"26",X"10",X"7D",X"9C",X"40",X"26",X"0B",X"8E",X"C9",X"21",X"86",
		X"00",X"BD",X"D0",X"55",X"7E",X"D0",X"0A",X"86",X"01",X"8E",X"C8",X"48",X"7E",X"F4",X"BE",X"8E",
		X"B4",X"12",X"10",X"8E",X"CA",X"A0",X"4F",X"B7",X"A1",X"77",X"B7",X"A1",X"76",X"A6",X"A4",X"44",
		X"44",X"44",X"44",X"8D",X"0C",X"A6",X"A0",X"84",X"0F",X"8D",X"06",X"10",X"8C",X"CC",X"0E",X"26",
		X"EC",X"85",X"0C",X"26",X"09",X"BB",X"A1",X"76",X"48",X"48",X"B7",X"A1",X"76",X"39",X"34",X"02",
		X"84",X"03",X"BB",X"A1",X"76",X"B7",X"A1",X"76",X"35",X"02",X"84",X"0C",X"44",X"44",X"CE",X"CC",
		X"0D",X"E6",X"C6",X"F7",X"A1",X"75",X"8C",X"B9",X"B2",X"25",X"04",X"30",X"89",X"FA",X"61",X"B6",
		X"A1",X"77",X"27",X"14",X"A6",X"84",X"84",X"F0",X"A7",X"84",X"B6",X"A1",X"75",X"84",X"0F",X"AA",
		X"84",X"A7",X"84",X"B6",X"A1",X"75",X"20",X"0D",X"73",X"A1",X"77",X"B6",X"A1",X"75",X"A7",X"84",
		X"7A",X"A1",X"76",X"2B",X"0B",X"30",X"88",X"18",X"7A",X"A1",X"76",X"2A",X"F1",X"7F",X"A1",X"77",
		X"7F",X"A1",X"76",X"39",X"D6",X"37",X"27",X"21",X"F1",X"A1",X"83",X"23",X"06",X"F7",X"A1",X"83",
		X"7C",X"A1",X"84",X"CE",X"C0",X"E9",X"8E",X"28",X"E5",X"BD",X"FF",X"CE",X"C0",X"02",X"02",X"4F",
		X"8E",X"48",X"E5",X"BD",X"FF",X"CE",X"C0",X"0E",X"02",X"86",X"10",X"8E",X"C8",X"F4",X"7E",X"F4",
		X"BE",X"86",X"FF",X"B7",X"A1",X"6A",X"86",X"02",X"8E",X"C9",X"2E",X"7E",X"F4",X"BE",X"86",X"0A",
		X"B7",X"A1",X"6A",X"7E",X"D0",X"0A",X"96",X"8C",X"27",X"06",X"BD",X"D3",X"DB",X"4A",X"20",X"F8",
		X"39",X"FE",X"74",X"40",X"11",X"11",X"85",X"81",X"81",X"81",X"88",X"82",X"82",X"22",X"24",X"22",
		X"42",X"24",X"24",X"24",X"44",X"24",X"44",X"49",X"44",X"94",X"41",X"88",X"14",X"41",X"88",X"14",
		X"41",X"88",X"94",X"41",X"88",X"94",X"49",X"88",X"14",X"98",X"58",X"94",X"98",X"18",X"94",X"46",
		X"66",X"62",X"42",X"42",X"42",X"42",X"25",X"24",X"24",X"68",X"24",X"24",X"24",X"26",X"11",X"18",
		X"18",X"58",X"18",X"58",X"81",X"44",X"98",X"81",X"44",X"98",X"81",X"44",X"98",X"14",X"94",X"94",
		X"16",X"22",X"24",X"24",X"A4",X"24",X"A4",X"24",X"24",X"24",X"24",X"24",X"FE",X"81",X"4A",X"42",
		X"42",X"42",X"42",X"44",X"99",X"99",X"41",X"88",X"14",X"41",X"88",X"14",X"46",X"24",X"24",X"24",
		X"24",X"24",X"24",X"A4",X"24",X"24",X"A4",X"22",X"42",X"4A",X"42",X"42",X"44",X"99",X"19",X"91",
		X"19",X"91",X"91",X"81",X"81",X"41",X"81",X"49",X"46",X"42",X"42",X"42",X"42",X"42",X"42",X"24",
		X"22",X"42",X"62",X"62",X"42",X"24",X"49",X"19",X"91",X"91",X"91",X"91",X"91",X"85",X"88",X"14",
		X"94",X"14",X"24",X"24",X"24",X"24",X"24",X"24",X"A4",X"24",X"24",X"41",X"81",X"81",X"18",X"18",
		X"94",X"41",X"88",X"14",X"14",X"24",X"42",X"24",X"24",X"24",X"24",X"24",X"24",X"24",X"44",X"98",
		X"18",X"18",X"18",X"58",X"89",X"44",X"18",X"85",X"14",X"24",X"14",X"24",X"A4",X"24",X"24",X"24",
		X"A4",X"24",X"28",X"24",X"44",X"18",X"19",X"19",X"81",X"41",X"81",X"14",X"24",X"24",X"24",X"24",
		X"22",X"42",X"42",X"64",X"41",X"85",X"81",X"81",X"18",X"19",X"41",X"89",X"44",X"42",X"22",X"42",
		X"24",X"24",X"24",X"24",X"24",X"44",X"18",X"14",X"98",X"11",X"81",X"81",X"41",X"89",X"44",X"42",
		X"22",X"42",X"24",X"24",X"24",X"24",X"24",X"44",X"18",X"94",X"41",X"88",X"89",X"44",X"49",X"88",
		X"14",X"41",X"88",X"14",X"14",X"24",X"24",X"24",X"26",X"62",X"66",X"26",X"24",X"18",X"91",X"91",
		X"19",X"18",X"14",X"18",X"14",X"14",X"24",X"14",X"2A",X"45",X"24",X"68",X"88",X"24",X"44",X"42",
		X"18",X"A8",X"82",X"44",X"A8",X"22",X"20",X"FE",X"87",X"40",X"44",X"11",X"88",X"24",X"FE",X"9A",
		X"3F",X"44",X"11",X"88",X"24",X"FE",X"C1",X"3F",X"44",X"44",X"44",X"11",X"11",X"11",X"11",X"88",
		X"88",X"88",X"22",X"22",X"22",X"20",X"FE",X"C3",X"45",X"22",X"22",X"44",X"11",X"81",X"50",X"FD",
		X"10",X"D1",X"BD",X"29",X"C2",X"9C",X"29",X"CB",X"EA",X"C2",X"8C",X"29",X"C2",X"81",X"0D",X"10",
		X"C2",X"8D",X"29",X"C2",X"9C",X"29",X"CB",X"EA",X"42",X"94",X"29",X"42",X"81",X"0C",X"3F",X"29",
		X"C2",X"94",X"C2",X"9C",X"29",X"C1",X"8D",X"A4",X"29",X"42",X"94",X"29",X"3F",X"3E",X"29",X"42",
		X"A4",X"29",X"4C",X"29",X"C1",X"8D",X"A4",X"2A",X"42",X"94",X"29",X"3E",X"3D",X"B6",X"B4",X"A2",
		X"4A",X"17",X"CA",X"16",X"C1",X"9C",X"B4",X"A7",X"A4",X"B1",X"7A",X"7A",X"3D",X"3C",X"B6",X"B4",
		X"B1",X"71",X"81",X"6B",X"16",X"C1",X"AC",X"A4",X"B6",X"B4",X"A2",X"4A",X"6B",X"3C",X"2F",X"B6",
		X"B4",X"29",X"62",X"85",X"C2",X"85",X"C1",X"AC",X"A4",X"B6",X"B4",X"28",X"62",X"A2",X"F2",X"EB",
		X"61",X"84",X"29",X"62",X"8E",X"28",X"E2",X"A4",X"B7",X"B4",X"28",X"62",X"A2",X"E2",X"DB",X"7B",
		X"42",X"96",X"28",X"4E",X"28",X"E2",X"B4",X"B6",X"B4",X"29",X"62",X"92",X"E2",X"CB",X"7B",X"52",
		X"96",X"28",X"4E",X"28",X"EB",X"41",X"A4",X"B7",X"B4",X"28",X"62",X"92",X"E1",X"FB",X"7B",X"5B",
		X"24",X"B1",X"6D",X"18",X"14",X"EB",X"51",X"94",X"B7",X"B4",X"18",X"17",X"29",X"2D",X"1E",X"B1",
		X"4B",X"4B",X"25",X"B1",X"6D",X"B1",X"5E",X"B5",X"1A",X"4B",X"61",X"84",X"B2",X"4B",X"41",X"82",
		X"C1",X"DB",X"14",X"B5",X"18",X"17",X"18",X"16",X"D1",X"81",X"4E",X"B6",X"19",X"4B",X"61",X"84",
		X"18",X"24",X"B4",X"18",X"1F",X"1C",X"38",X"53",X"84",X"B1",X"6E",X"2B",X"CB",X"61",X"94",X"38",
		X"42",X"B4",X"18",X"41",X"81",X"EF",X"39",X"43",X"85",X"B1",X"6E",X"2B",X"CB",X"71",X"84",X"38",
		X"43",X"84",X"B6",X"18",X"1C",X"E3",X"95",X"38",X"41",X"81",X"6D",X"38",X"CB",X"C6",X"19",X"42",
		X"B5",X"38",X"4B",X"61",X"8F",X"D3",X"95",X"38",X"5B",X"51",X"F3",X"8C",X"BD",X"61",X"84",X"2A",
		X"63",X"85",X"B6",X"18",X"ED",X"38",X"53",X"94",X"18",X"51",X"F3",X"8C",X"BD",X"7B",X"42",X"91",
		X"42",X"B5",X"18",X"7B",X"DC",X"21",X"51",X"F3",X"4C",X"7E",X"30",X"6C",X"C2",X"14",X"2C",X"34",
		X"C7",X"E1",X"07",X"C1",X"35",X"CC",X"21",X"42",X"C3",X"4C",X"7F",X"10",X"6C",X"13",X"5C",X"C1",
		X"35",X"C1",X"52",X"C3",X"4C",X"7F",X"15",X"C2",X"7D",X"34",X"C1",X"5C",X"17",X"CC",X"36",X"C3",
		X"5C",X"14",X"2D",X"34",X"C7",X"1C",X"14",X"C2",X"6E",X"34",X"D1",X"4E",X"15",X"CC",X"36",X"C3",
		X"5C",X"14",X"2D",X"34",X"C7",X"1C",X"14",X"C2",X"51",X"C2",X"7D",X"14",X"F1",X"4C",X"22",X"CC",
		X"00",X"3E",X"41",X"41",X"22",X"00",X"3E",X"41",X"41",X"3E",X"00",X"7F",X"09",X"09",X"06",X"00",
		X"03",X"04",X"78",X"04",X"03",X"00",X"7F",X"09",X"19",X"66",X"00",X"41",X"7F",X"41",X"00",X"3E",
		X"41",X"49",X"3A",X"00",X"7F",X"08",X"08",X"7F",X"00",X"01",X"01",X"7F",X"01",X"01",X"00",X"1C",
		X"22",X"5D",X"63",X"55",X"22",X"1C",X"22",X"7F",X"4B",X"45",X"22",X"1C",X"00",X"00",X"00",X"42",
		X"7F",X"40",X"00",X"26",X"49",X"49",X"3E",X"00",X"36",X"49",X"49",X"36",X"00",X"3E",X"41",X"41",
		X"3E",X"43",X"30",X"1C",X"70",X"3C",X"70",X"5F",X"70",X"1C",X"A8",X"40",X"A8",X"5C",X"A8",X"C0",
		X"EB",X"C0",X"DD",X"C0",X"DF",X"C0",X"E7",X"C0",X"E3",X"C0",X"E1",X"C0",X"E5",X"60",X"00",X"60",
		X"00",X"62",X"00",X"98",X"00",X"98",X"00",X"9A",X"00",X"F9",X"85",X"F8",X"CE",X"F9",X"A3",X"F9",
		X"29",X"F8",X"F7",X"F9",X"7B",X"09",X"00",X"11",X"00",X"19",X"80",X"09",X"60",X"11",X"60",X"19",
		X"E0",X"44",X"33",X"CC",X"33",X"33",X"33",X"88",X"88",X"CC",X"CC",X"24",X"24",X"CE",X"00",X"00",
		X"C6",X"08",X"8E",X"B0",X"5D",X"EF",X"94",X"EF",X"98",X"02",X"EF",X"98",X"04",X"EF",X"98",X"06",
		X"3A",X"9C",X"97",X"25",X"F0",X"AE",X"9F",X"A0",X"97",X"27",X"08",X"EF",X"84",X"6F",X"02",X"EF",
		X"89",X"FF",X"00",X"DC",X"20",X"83",X"6D",X"40",X"DD",X"73",X"44",X"44",X"CE",X"CD",X"69",X"C6",
		X"03",X"3D",X"33",X"CB",X"96",X"BA",X"85",X"02",X"26",X"22",X"86",X"30",X"10",X"8E",X"B1",X"25",
		X"8E",X"00",X"00",X"AF",X"B4",X"37",X"14",X"ED",X"A4",X"AF",X"B1",X"4C",X"8E",X"00",X"00",X"AF",
		X"B4",X"37",X"14",X"ED",X"A4",X"AF",X"B1",X"4C",X"81",X"70",X"26",X"E4",X"8E",X"4C",X"09",X"CC",
		X"90",X"90",X"ED",X"84",X"ED",X"88",X"1D",X"8E",X"53",X"09",X"CC",X"09",X"09",X"ED",X"84",X"ED",
		X"88",X"1D",X"8E",X"A0",X"65",X"CE",X"B0",X"5D",X"8D",X"3A",X"8E",X"A0",X"6B",X"8D",X"35",X"DF",
		X"97",X"DC",X"BF",X"44",X"44",X"44",X"44",X"54",X"54",X"54",X"C3",X"4B",X"07",X"ED",X"C4",X"AE",
		X"C4",X"CC",X"90",X"99",X"ED",X"84",X"A7",X"02",X"86",X"09",X"A7",X"89",X"FF",X"01",X"39",X"EC",
		X"0A",X"93",X"73",X"44",X"44",X"E6",X"0C",X"54",X"54",X"54",X"C3",X"30",X"07",X"ED",X"C4",X"EC",
		X"88",X"12",X"ED",X"D1",X"AE",X"84",X"26",X"E7",X"39",X"25",X"70",X"07",X"26",X"77",X"00",X"26",
		X"07",X"70",X"24",X"07",X"70",X"23",X"07",X"70",X"23",X"70",X"07",X"24",X"07",X"70",X"25",X"70",
		X"07",X"26",X"77",X"00",X"25",X"07",X"70",X"24",X"07",X"70",X"23",X"07",X"70",X"21",X"07",X"70",
		X"22",X"70",X"07",X"24",X"77",X"00",X"24",X"70",X"07",X"26",X"77",X"00",X"26",X"77",X"00",X"25",
		X"77",X"00",X"25",X"70",X"07",X"26",X"77",X"00",X"24",X"07",X"70",X"23",X"70",X"07",X"25",X"77",
		X"00",X"26",X"70",X"07",X"26",X"77",X"00",X"26",X"77",X"00",X"25",X"07",X"70",X"23",X"07",X"70",
		X"22",X"07",X"70",X"21",X"77",X"00",X"21",X"70",X"07",X"23",X"70",X"07",X"25",X"70",X"07",X"25",
		X"07",X"70",X"25",X"77",X"00",X"25",X"77",X"00",X"24",X"77",X"00",X"22",X"07",X"70",X"20",X"07",
		X"70",X"1E",X"07",X"70",X"1C",X"07",X"70",X"1D",X"70",X"07",X"1F",X"70",X"07",X"21",X"70",X"07",
		X"22",X"70",X"07",X"24",X"70",X"07",X"26",X"70",X"07",X"26",X"77",X"00",X"26",X"77",X"00",X"26",
		X"77",X"00",X"26",X"77",X"00",X"26",X"77",X"00",X"25",X"77",X"00",X"25",X"70",X"07",X"26",X"77",
		X"00",X"24",X"07",X"70",X"23",X"77",X"00",X"24",X"77",X"00",X"22",X"07",X"70",X"23",X"70",X"07",
		X"22",X"07",X"70",X"21",X"70",X"07",X"23",X"70",X"07",X"25",X"70",X"07",X"26",X"77",X"00",X"26",
		X"07",X"70",X"24",X"07",X"70",X"23",X"07",X"70",X"23",X"70",X"07",X"24",X"07",X"70",X"25",X"70",
		X"07",X"26",X"77",X"00",X"25",X"07",X"70",X"24",X"07",X"70",X"23",X"07",X"70",X"21",X"07",X"70",
		X"22",X"70",X"07",X"24",X"77",X"00",X"24",X"70",X"07",X"26",X"77",X"00",X"26",X"77",X"00",X"25",
		X"77",X"00",X"25",X"70",X"07",X"26",X"77",X"00",X"24",X"07",X"70",X"23",X"70",X"07",X"25",X"77",
		X"00",X"26",X"70",X"07",X"26",X"77",X"00",X"26",X"77",X"00",X"25",X"07",X"70",X"23",X"07",X"70",
		X"22",X"07",X"70",X"21",X"77",X"00",X"21",X"70",X"07",X"23",X"70",X"07",X"25",X"70",X"07",X"25",
		X"07",X"70",X"25",X"77",X"00",X"25",X"77",X"00",X"24",X"77",X"00",X"22",X"07",X"70",X"20",X"07",
		X"70",X"1E",X"07",X"70",X"1C",X"07",X"70",X"1D",X"70",X"07",X"1F",X"70",X"07",X"21",X"70",X"07",
		X"22",X"70",X"07",X"24",X"70",X"07",X"26",X"70",X"07",X"26",X"77",X"00",X"26",X"77",X"00",X"26",
		X"77",X"00",X"26",X"77",X"00",X"26",X"77",X"00",X"25",X"77",X"00",X"25",X"70",X"07",X"26",X"77",
		X"00",X"24",X"07",X"70",X"23",X"77",X"00",X"24",X"77",X"00",X"22",X"07",X"70",X"23",X"70",X"07",
		X"22",X"07",X"70",X"21",X"70",X"07",X"23",X"70",X"07",X"80",X"00",X"00",X"30",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"00",X"FE",
		X"C3",X"00",X"00",X"00",X"00",X"D6",X"66",X"00",X"00",X"00",X"00",X"66",X"66",X"39",X"00",X"06",
		X"66",X"66",X"88",X"68",X"66",X"66",X"66",X"88",X"88",X"88",X"00",X"60",X"63",X"30",X"63",X"00",
		X"06",X"26",X"68",X"28",X"60",X"66",X"66",X"86",X"00",X"00",X"66",X"66",X"00",X"00",X"ED",X"66",
		X"00",X"00",X"00",X"63",X"90",X"09",X"90",X"99",X"99",X"99",X"90",X"CC",X"90",X"11",X"00",X"11",
		X"10",X"11",X"00",X"10",X"10",X"10",X"00",X"10",X"00",X"11",X"10",X"11",X"00",X"11",X"00",X"10",
		X"00",X"10",X"10",X"10",X"00",X"11",X"10",X"10",X"10",X"11",X"00",X"10",X"10",X"10",X"10",X"10",
		X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"11",X"01",X"11",X"00",X"11",X"00",X"01",X"01",X"01",
		X"00",X"01",X"00",X"11",X"00",X"11",X"01",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"11",
		X"01",X"01",X"01",X"11",X"00",X"FF",X"F0",X"FF",X"00",X"FF",X"00",X"F0",X"00",X"F0",X"F0",X"F0",
		X"00",X"EE",X"E0",X"E0",X"E0",X"EE",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"DD",X"D0",X"D0",
		X"D0",X"DD",X"00",X"D0",X"D0",X"D0",X"D0",X"D0",X"00",X"0F",X"0F",X"0F",X"00",X"0F",X"00",X"FF",
		X"00",X"FF",X"0F",X"FF",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"EE",X"0E",X"0E",X"0E",X"EE",
		X"00",X"0D",X"0D",X"0D",X"0D",X"0D",X"00",X"DD",X"0D",X"0D",X"0D",X"DD",X"00",X"1C",X"0D",X"7F",
		X"E7",X"70",X"00",X"0F",X"71",X"71",X"07",X"DC",X"77",X"7C",X"0D",X"71",X"C7",X"77",X"DE",X"07",
		X"71",X"17",X"17",X"DE",X"F7",X"71",X"17",X"71",X"7C",X"DE",X"F0",X"07",X"77",X"C7",X"71",X"17",
		X"70",X"70",X"7C",X"D7",X"77",X"77",X"70",X"01",X"CD",X"FF",X"D7",X"70",X"F0",X"00",X"00",X"00",
		X"C5",X"FB",X"7E",X"CA",X"A7",X"7E",X"CA",X"B2",X"7E",X"CA",X"BD",X"7E",X"CA",X"C8",X"7E",X"CB",
		X"C1",X"7E",X"CB",X"CC",X"7E",X"CB",X"D7",X"7E",X"CB",X"E2",X"7E",X"CA",X"79",X"7E",X"CA",X"81",
		X"7E",X"CA",X"51",X"7E",X"CA",X"58",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5B",
		X"FF",X"C0",X"BD",X"C0",X"BF",X"C0",X"C1",X"00",X"00",X"C0",X"C1",X"00",X"00",X"C0",X"C3",X"00",
		X"00",X"C0",X"C5",X"00",X"00",X"C0",X"C5",X"00",X"00",X"C0",X"C7",X"00",X"00",X"C0",X"C3",X"00",
		X"00",X"C0",X"C9",X"00",X"00",X"C0",X"CB",X"C0",X"CD",X"C0",X"CF",X"00",X"00",X"C0",X"BD",X"C0",
		X"D1",X"C0",X"D3",X"C0",X"D5",X"C0",X"DB",X"00",X"00",X"C1",X"07",X"C1",X"0D",X"C1",X"11",X"C1",
		X"13",X"C1",X"15",X"C1",X"19",X"C1",X"1D",X"C1",X"21",X"C1",X"27",X"C1",X"2B",X"C1",X"33",X"C1",
		X"4D",X"C1",X"53",X"C1",X"6D",X"C1",X"88",X"C1",X"92",X"C1",X"96",X"C1",X"9C",X"C1",X"A0",X"C1",
		X"A2",X"C1",X"A6",X"C1",X"A8",X"C1",X"AC",X"C1",X"B0",X"C1",X"B2",X"C1",X"B4",X"C1",X"B6",X"C1",
		X"B8",X"C1",X"BC",X"C1",X"BE",X"C1",X"C2",X"C1",X"C6",X"C1",X"C8",X"C1",X"CA",X"C1",X"CC",X"C1",
		X"CE",X"C1",X"D0",X"C1",X"D2",X"C1",X"D4",X"C1",X"D6",X"C1",X"D8",X"C1",X"DA",X"C1",X"EA",X"C1",
		X"F8",X"C2",X"00",X"C2",X"08",X"C2",X"10",X"C2",X"1A",X"C2",X"24",X"C2",X"2C",X"C2",X"34",X"C2",
		X"3E",X"C2",X"48",X"C2",X"52",X"C2",X"5A",X"C2",X"64",X"C2",X"68",X"C2",X"74",X"C2",X"7E",X"C2",
		X"85",X"C2",X"8C",X"C2",X"93",X"C2",X"9A",X"C2",X"A1",X"C2",X"A8",X"C2",X"AA",X"C2",X"AC",X"C2",
		X"B4",X"C2",X"B8",X"C2",X"BC",X"C2",X"BE",X"C2",X"C6",X"C2",X"D2",X"C2",X"D6",X"C2",X"D8",X"C3",
		X"01",X"C3",X"0B",X"C3",X"21",X"C3",X"2B",X"C4",X"64",X"C5",X"8D",X"C4",X"50",X"C5",X"BB",X"C4",
		X"D1",X"C5",X"2D",X"C5",X"1B",X"C5",X"2D",X"C4",X"04",X"C5",X"1B",X"C4",X"04",X"C4",X"15",X"C4",
		X"E0",X"C3",X"3E",X"C5",X"31",X"C4",X"D1",X"C5",X"1B",X"C5",X"81",X"C4",X"CA",X"C5",X"1B",X"C3",
		X"F8",X"C3",X"C6",X"C3",X"93",X"C5",X"1B",X"C4",X"04",X"06",X"28",X"A0",X"C5",X"81",X"C4",X"AD",
		X"C3",X"66",X"C3",X"F0",X"07",X"C5",X"DA",X"C3",X"98",X"C3",X"CF",X"C4",X"D8",X"C3",X"93",X"C5",
		X"1B",X"C4",X"D1",X"C4",X"A4",X"C5",X"1B",X"C4",X"04",X"03",X"FE",X"C3",X"81",X"04",X"10",X"02",
		X"F8",X"C3",X"93",X"C5",X"1B",X"C3",X"7D",X"C4",X"CD",X"C3",X"66",X"C5",X"86",X"C3",X"9D",X"C5",
		X"1B",X"C5",X"81",X"04",X"30",X"02",X"E8",X"C5",X"C3",X"C3",X"9D",X"C3",X"61",X"C4",X"50",X"07",
		X"03",X"FC",X"C3",X"9D",X"C5",X"1B",X"C4",X"04",X"C3",X"49",X"C5",X"81",X"07",X"07",X"03",X"04",
		X"C5",X"54",X"C5",X"7A",X"C5",X"81",X"C4",X"9C",X"C5",X"81",X"C4",X"E5",X"C3",X"55",X"C5",X"C0",
		X"C3",X"36",X"C5",X"27",X"C3",X"98",X"C4",X"35",X"C4",X"8B",X"C3",X"98",X"C3",X"85",X"C3",X"98",
		X"C4",X"75",X"C4",X"75",X"C4",X"0C",X"C5",X"9C",X"C5",X"4E",X"C3",X"69",X"C4",X"45",X"C5",X"B7",
		X"C4",X"F5",X"C4",X"D4",X"C4",X"EE",X"C5",X"1F",X"C3",X"D4",X"C5",X"C0",X"C4",X"75",X"C4",X"75",
		X"C4",X"75",X"C4",X"75",X"C4",X"75",X"C4",X"75",X"C4",X"75",X"C5",X"0B",X"C3",X"36",X"C5",X"DA",
		X"C5",X"7A",X"C5",X"45",X"C4",X"11",X"03",X"FE",X"C3",X"83",X"C3",X"55",X"C4",X"11",X"C3",X"4F",
		X"03",X"FE",X"C3",X"81",X"C4",X"15",X"C3",X"2B",X"C4",X"95",X"C4",X"11",X"C5",X"2D",X"C5",X"81",
		X"C3",X"55",X"C4",X"11",X"C5",X"1B",X"C5",X"81",X"C3",X"55",X"C5",X"AD",X"C3",X"FF",X"C5",X"81",
		X"C3",X"55",X"C4",X"11",X"C3",X"93",X"C5",X"1B",X"C5",X"81",X"C3",X"55",X"C4",X"11",X"C3",X"9D",
		X"C5",X"1B",X"C5",X"81",X"C3",X"55",X"C4",X"11",X"C3",X"49",X"C5",X"81",X"C3",X"55",X"C4",X"11",
		X"C5",X"7A",X"C5",X"81",X"C4",X"95",X"C5",X"AD",X"C5",X"81",X"C4",X"59",X"C5",X"5A",X"C3",X"55",
		X"C4",X"11",X"C4",X"9C",X"C5",X"81",X"C4",X"E5",X"C4",X"95",X"C5",X"AD",X"C5",X"67",X"C5",X"97",
		X"C4",X"E5",X"C3",X"55",X"C4",X"11",X"C4",X"15",X"C4",X"E0",X"C4",X"95",X"C5",X"AD",X"C5",X"67",
		X"C5",X"97",X"C3",X"2B",X"C5",X"D1",X"C3",X"BD",X"C5",X"0B",X"C3",X"36",X"C5",X"AD",X"C5",X"67",
		X"C5",X"97",X"C5",X"81",X"C5",X"0B",X"C4",X"35",X"C5",X"AD",X"C4",X"90",X"C3",X"8C",X"C4",X"84",
		X"07",X"03",X"06",X"C4",X"B9",X"C4",X"B2",X"07",X"03",X"06",X"C4",X"B9",X"C4",X"FD",X"07",X"03",
		X"00",X"C4",X"C5",X"C3",X"6E",X"07",X"03",X"06",X"C4",X"C1",X"C5",X"72",X"07",X"03",X"08",X"C4",
		X"B9",X"C3",X"5A",X"07",X"03",X"06",X"C4",X"BD",X"C3",X"B4",X"C5",X"36",X"C3",X"D9",X"07",X"07",
		X"03",X"0C",X"C5",X"02",X"C4",X"EE",X"C4",X"D4",X"C4",X"EE",X"C5",X"B7",X"C3",X"75",X"C5",X"0B",
		X"C4",X"D4",X"C4",X"EE",X"C5",X"61",X"C5",X"0B",X"C4",X"D4",X"C4",X"DD",X"C5",X"B7",X"C4",X"EE",
		X"C5",X"61",X"C3",X"42",X"C5",X"CC",X"C3",X"A3",X"C5",X"DF",X"C4",X"30",X"C5",X"11",X"C4",X"11",
		X"07",X"C5",X"93",X"C3",X"BD",X"C4",X"23",X"07",X"07",X"C5",X"3E",X"C4",X"6C",X"C5",X"DA",X"C5",
		X"C0",X"C3",X"D4",X"C5",X"6C",X"07",X"07",X"C5",X"0B",X"C4",X"0C",X"C5",X"AD",X"C3",X"EA",X"C4",
		X"64",X"A0",X"00",X"02",X"08",X"A0",X"02",X"02",X"10",X"A0",X"04",X"C4",X"23",X"06",X"22",X"68",
		X"C5",X"B0",X"02",X"3E",X"C3",X"3E",X"C5",X"A8",X"07",X"03",X"FC",X"C4",X"1A",X"02",X"3D",X"C4",
		X"1A",X"A0",X"06",X"02",X"05",X"A0",X"08",X"02",X"13",X"A0",X"0C",X"41",X"44",X"4A",X"55",X"53",
		X"54",X"4D",X"45",X"4E",X"54",X"2F",X"41",X"44",X"56",X"41",X"4E",X"43",X"45",X"2F",X"41",X"4C",
		X"4C",X"2F",X"41",X"54",X"54",X"41",X"43",X"4B",X"2F",X"41",X"55",X"44",X"49",X"4F",X"2F",X"41",
		X"55",X"44",X"49",X"54",X"2F",X"41",X"55",X"54",X"4F",X"2F",X"42",X"41",X"49",X"54",X"45",X"52",
		X"2F",X"42",X"41",X"52",X"53",X"2F",X"42",X"45",X"2F",X"42",X"4F",X"4D",X"42",X"2F",X"42",X"4F",
		X"4D",X"42",X"45",X"52",X"2F",X"42",X"4F",X"4E",X"55",X"53",X"20",X"58",X"2F",X"43",X"41",X"4E",
		X"2F",X"2C",X"2F",X"3A",X"2F",X"43",X"45",X"4E",X"54",X"45",X"52",X"2F",X"43",X"48",X"41",X"4E",
		X"47",X"45",X"2F",X"43",X"4D",X"4F",X"53",X"2F",X"43",X"4F",X"49",X"4E",X"2F",X"43",X"4F",X"4C",
		X"4F",X"52",X"2F",X"43",X"4F",X"4D",X"50",X"4C",X"45",X"54",X"45",X"44",X"2F",X"43",X"52",X"45",
		X"44",X"49",X"54",X"2F",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"3A",X"2F",X"44",X"45",X"46",
		X"45",X"4E",X"44",X"45",X"52",X"2F",X"44",X"45",X"54",X"45",X"43",X"54",X"45",X"44",X"2F",X"44",
		X"4F",X"4F",X"52",X"2F",X"44",X"4F",X"57",X"4E",X"2F",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",
		X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"2F",X"45",X"4E",X"54",X"45",X"52",X"2F",
		X"45",X"4E",X"54",X"45",X"52",X"45",X"44",X"2F",X"45",X"52",X"52",X"4F",X"52",X"53",X"2F",X"45",
		X"58",X"49",X"54",X"2F",X"46",X"41",X"49",X"4C",X"55",X"52",X"45",X"2F",X"46",X"49",X"52",X"45",
		X"2F",X"46",X"4F",X"52",X"2F",X"47",X"41",X"4D",X"45",X"2F",X"47",X"52",X"45",X"41",X"54",X"45",
		X"53",X"54",X"2F",X"48",X"41",X"4C",X"4C",X"20",X"4F",X"46",X"20",X"46",X"41",X"4D",X"45",X"2F",
		X"48",X"41",X"56",X"45",X"2F",X"48",X"49",X"47",X"48",X"53",X"43",X"4F",X"52",X"45",X"20",X"52",
		X"45",X"53",X"45",X"54",X"2F",X"48",X"59",X"50",X"45",X"52",X"53",X"50",X"41",X"43",X"45",X"2F",
		X"49",X"4E",X"44",X"49",X"43",X"41",X"54",X"45",X"2F",X"49",X"4E",X"44",X"49",X"56",X"49",X"44",
		X"55",X"41",X"4C",X"2F",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"2F",X"49",X"4E",X"49",X"54",
		X"49",X"41",X"4C",X"53",X"2F",X"49",X"4E",X"56",X"41",X"4C",X"49",X"44",X"20",X"53",X"57",X"49",
		X"54",X"43",X"48",X"2F",X"4C",X"41",X"4E",X"44",X"45",X"52",X"2F",X"4C",X"45",X"46",X"54",X"2F",
		X"4D",X"41",X"4B",X"45",X"2F",X"4D",X"41",X"4E",X"55",X"41",X"4C",X"2F",X"4D",X"4F",X"4E",X"49",
		X"54",X"4F",X"52",X"2F",X"4D",X"55",X"4C",X"54",X"49",X"50",X"4C",X"45",X"2F",X"4D",X"55",X"53",
		X"54",X"2F",X"4D",X"55",X"54",X"41",X"4E",X"54",X"2F",X"31",X"35",X"30",X"2F",X"32",X"30",X"30",
		X"2F",X"32",X"35",X"30",X"2F",X"31",X"30",X"30",X"30",X"2F",X"4E",X"4F",X"2F",X"4E",X"4F",X"54",
		X"2F",X"4F",X"4B",X"2F",X"4F",X"4E",X"45",X"2F",X"4F",X"50",X"45",X"4E",X"2F",X"4F",X"52",X"2F",
		X"4F",X"56",X"45",X"52",X"2F",X"50",X"41",X"54",X"54",X"45",X"52",X"4E",X"53",X"2F",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"2F",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"2F",X"20",X"50",X"4F",
		X"44",X"2F",X"50",X"52",X"45",X"53",X"45",X"4E",X"54",X"53",X"2F",X"50",X"52",X"45",X"53",X"53",
		X"2F",X"51",X"55",X"41",X"4C",X"49",X"46",X"49",X"45",X"44",X"2F",X"52",X"41",X"4D",X"2F",X"52",
		X"45",X"56",X"45",X"52",X"53",X"45",X"2F",X"52",X"49",X"47",X"48",X"54",X"2F",X"52",X"4F",X"4D",
		X"2F",X"52",X"4F",X"4D",X"53",X"2F",X"53",X"43",X"41",X"4E",X"4E",X"45",X"52",X"2F",X"53",X"45",
		X"4C",X"45",X"43",X"54",X"2F",X"53",X"45",X"54",X"2F",X"53",X"4C",X"41",X"4D",X"2F",X"53",X"4D",
		X"41",X"52",X"54",X"2F",X"53",X"4F",X"55",X"4E",X"44",X"2F",X"53",X"4F",X"55",X"4E",X"44",X"53",
		X"2F",X"53",X"54",X"41",X"52",X"54",X"2F",X"53",X"54",X"45",X"50",X"2F",X"53",X"54",X"49",X"43",
		X"4B",X"2F",X"53",X"57",X"41",X"52",X"4D",X"45",X"52",X"2F",X"53",X"57",X"49",X"54",X"43",X"48",
		X"2F",X"54",X"45",X"53",X"54",X"2F",X"54",X"45",X"53",X"54",X"45",X"44",X"2F",X"54",X"45",X"53",
		X"54",X"53",X"2F",X"54",X"48",X"45",X"2F",X"54",X"48",X"52",X"55",X"2F",X"54",X"48",X"52",X"55",
		X"53",X"54",X"2F",X"54",X"49",X"4C",X"54",X"2F",X"54",X"49",X"4D",X"45",X"2F",X"54",X"4F",X"2F",
		X"54",X"4F",X"44",X"41",X"59",X"53",X"2F",X"54",X"57",X"4F",X"2F",X"55",X"4E",X"49",X"54",X"2F",
		X"55",X"50",X"2F",X"56",X"45",X"52",X"54",X"49",X"43",X"41",X"4C",X"2F",X"57",X"41",X"56",X"45",
		X"2F",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"2F",X"57",X"49",X"54",X"48",X"2F",X"59",
		X"4F",X"55",X"2F",X"01",X"08",X"C6",X"97",X"01",X"08",X"C6",X"AF",X"01",X"08",X"C6",X"B7",X"03",
		X"08",X"C7",X"BF",X"01",X"08",X"C6",X"BF",X"03",X"08",X"C7",X"BF",X"03",X"08",X"C6",X"C7",X"03",
		X"08",X"C6",X"DF",X"03",X"08",X"C6",X"F7",X"03",X"08",X"C7",X"0F",X"03",X"08",X"C7",X"27",X"03",
		X"08",X"C7",X"3F",X"03",X"08",X"C7",X"57",X"03",X"08",X"C7",X"6F",X"03",X"08",X"C7",X"87",X"03",
		X"08",X"C7",X"9F",X"01",X"08",X"C7",X"B7",X"03",X"08",X"C7",X"BF",X"03",X"08",X"C6",X"97",X"03",
		X"08",X"C7",X"D7",X"03",X"08",X"C7",X"EF",X"03",X"08",X"C8",X"07",X"03",X"08",X"C8",X"1F",X"03",
		X"08",X"C8",X"37",X"03",X"08",X"C8",X"4F",X"03",X"08",X"C8",X"67",X"03",X"08",X"C8",X"7F",X"02",
		X"08",X"C8",X"97",X"03",X"08",X"C8",X"A7",X"03",X"08",X"C8",X"BF",X"03",X"08",X"C8",X"D7",X"04",
		X"08",X"C8",X"EF",X"03",X"08",X"C9",X"0F",X"03",X"08",X"C9",X"27",X"03",X"08",X"C9",X"3F",X"03",
		X"08",X"C9",X"57",X"03",X"08",X"C9",X"6F",X"03",X"08",X"C9",X"87",X"03",X"08",X"C9",X"9F",X"03",
		X"08",X"C9",X"B7",X"03",X"08",X"C9",X"CF",X"04",X"08",X"C9",X"E7",X"03",X"08",X"CA",X"07",X"03",
		X"08",X"CA",X"1F",X"03",X"08",X"CA",X"37",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"01",X"01",X"01",X"01",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"10",X"00",X"00",X"00",X"00",X"00",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"00",X"11",
		X"00",X"00",X"01",X"10",X"00",X"11",X"00",X"11",X"11",X"11",X"10",X"00",X"00",X"11",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"01",
		X"10",X"00",X"11",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"01",
		X"01",X"01",X"01",X"00",X"00",X"01",X"00",X"11",X"10",X"10",X"11",X"00",X"00",X"11",X"00",X"11",
		X"00",X"00",X"11",X"01",X"01",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",
		X"10",X"10",X"11",X"10",X"10",X"11",X"00",X"11",X"00",X"00",X"11",X"01",X"01",X"11",X"00",X"01",
		X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"11",X"00",X"00",X"01",X"11",X"10",X"10",X"00",X"11",
		X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"00",X"11",
		X"10",X"10",X"11",X"10",X"10",X"11",X"00",X"11",X"01",X"01",X"10",X"01",X"01",X"11",X"00",X"01",
		X"01",X"01",X"01",X"00",X"00",X"01",X"00",X"11",X"10",X"10",X"11",X"00",X"00",X"11",X"00",X"11",
		X"01",X"01",X"11",X"01",X"01",X"11",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"01",X"01",X"00",X"01",X"00",X"11",
		X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",
		X"10",X"10",X"10",X"10",X"10",X"11",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"10",
		X"11",X"11",X"11",X"11",X"11",X"10",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",
		X"10",X"10",X"11",X"10",X"10",X"11",X"00",X"11",X"00",X"00",X"10",X"00",X"00",X"11",X"00",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"10",X"10",X"11",X"10",X"10",X"10",X"00",X"11",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",
		X"10",X"10",X"10",X"10",X"10",X"11",X"00",X"11",X"00",X"00",X"11",X"01",X"01",X"11",X"00",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"10",X"10",X"10",X"11",X"10",X"10",X"10",X"00",X"01",
		X"01",X"01",X"11",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"01",X"11",X"01",X"00",X"00",X"00",X"01",
		X"10",X"00",X"00",X"00",X"10",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"10",
		X"10",X"10",X"10",X"10",X"10",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"11",
		X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"11",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",
		X"10",X"10",X"10",X"10",X"10",X"11",X"00",X"11",X"01",X"01",X"01",X"01",X"01",X"11",X"00",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"10",X"10",X"11",X"10",X"10",X"10",X"00",X"11",
		X"01",X"01",X"11",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",
		X"10",X"10",X"10",X"10",X"10",X"11",X"00",X"11",X"01",X"01",X"01",X"01",X"11",X"11",X"10",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"11",X"10",X"10",X"11",X"10",X"10",X"10",X"00",X"11",
		X"01",X"01",X"11",X"10",X"01",X"01",X"00",X"01",X"01",X"01",X"01",X"00",X"00",X"01",X"00",X"11",
		X"10",X"10",X"11",X"00",X"00",X"11",X"00",X"11",X"00",X"00",X"11",X"11",X"11",X"11",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"10",
		X"10",X"10",X"10",X"10",X"10",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"11",X"00",X"01",
		X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"00",X"01",
		X"01",X"01",X"01",X"01",X"10",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"10",
		X"10",X"10",X"10",X"10",X"10",X"01",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"01",X"00",X"10",
		X"10",X"10",X"10",X"10",X"10",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"00",X"10",X"01",X"10",X"00",X"00",X"00",X"01",X"01",X"10",X"00",X"10",X"01",X"01",X"00",X"01",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"01",X"01",X"01",X"00",X"01",
		X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"01",X"01",X"00",X"11",
		X"00",X"01",X"10",X"00",X"00",X"11",X"00",X"11",X"10",X"00",X"00",X"00",X"00",X"11",X"00",X"84",
		X"FF",X"34",X"70",X"CE",X"C0",X"D9",X"20",X"05",X"34",X"70",X"CE",X"C0",X"BB",X"8E",X"18",X"CE",
		X"BD",X"CA",X"A7",X"EE",X"A1",X"27",X"06",X"8E",X"10",X"DA",X"BD",X"CA",X"A7",X"EE",X"A1",X"27",
		X"06",X"8E",X"10",X"E4",X"BD",X"CA",X"A7",X"35",X"F0",X"34",X"77",X"10",X"8E",X"FF",X"B6",X"20",
		X"06",X"34",X"77",X"10",X"8E",X"FF",X"B3",X"CC",X"CA",X"ED",X"10",X"9F",X"3D",X"DD",X"3F",X"9F",
		X"50",X"9F",X"4E",X"8E",X"01",X"0A",X"9F",X"4C",X"0F",X"58",X"EE",X"65",X"DF",X"54",X"33",X"C8",
		X"20",X"DF",X"56",X"DF",X"52",X"20",X"46",X"34",X"77",X"10",X"8E",X"FF",X"B3",X"CC",X"CA",X"ED",
		X"20",X"1F",X"34",X"77",X"10",X"8E",X"FF",X"B6",X"CC",X"CA",X"ED",X"20",X"14",X"34",X"77",X"10",
		X"8E",X"FF",X"B3",X"CC",X"CB",X"5F",X"20",X"09",X"34",X"77",X"10",X"8E",X"FF",X"B6",X"CC",X"CB",
		X"5F",X"10",X"9F",X"3D",X"DD",X"3F",X"0D",X"52",X"26",X"13",X"9F",X"50",X"9F",X"4E",X"8E",X"01",
		X"0A",X"9F",X"4C",X"0F",X"58",X"AE",X"42",X"9F",X"56",X"AE",X"C4",X"20",X"21",X"0D",X"58",X"26",
		X"0E",X"9E",X"54",X"E6",X"80",X"C1",X"2F",X"26",X"30",X"C6",X"20",X"D7",X"58",X"20",X"2A",X"0F",
		X"58",X"9E",X"52",X"9C",X"56",X"26",X"07",X"0F",X"52",X"35",X"77",X"1A",X"01",X"39",X"EE",X"81",
		X"2B",X"11",X"30",X"1F",X"1F",X"30",X"81",X"08",X"22",X"ED",X"48",X"10",X"8E",X"CB",X"64",X"AD",
		X"B6",X"20",X"E0",X"9F",X"52",X"DF",X"54",X"20",X"C4",X"9F",X"54",X"C0",X"20",X"C1",X"01",X"23",
		X"16",X"C1",X"0B",X"23",X"10",X"C0",X"0A",X"C1",X"10",X"23",X"0C",X"C1",X"14",X"23",X"06",X"C0",
		X"04",X"C1",X"2C",X"23",X"02",X"C6",X"03",X"58",X"58",X"8E",X"C5",X"E3",X"3A",X"1F",X"12",X"DC",
		X"50",X"9E",X"3D",X"AD",X"84",X"AB",X"A4",X"9B",X"4C",X"97",X"50",X"9E",X"3F",X"6E",X"84",X"35",
		X"77",X"1C",X"FE",X"39",X"CB",X"76",X"CB",X"7B",X"CB",X"80",X"CB",X"87",X"CB",X"8E",X"CB",X"95",
		X"CB",X"9C",X"CB",X"A3",X"CB",X"AC",X"A6",X"80",X"97",X"4C",X"39",X"E6",X"80",X"D7",X"4D",X"39",
		X"96",X"4E",X"AB",X"80",X"97",X"50",X"39",X"96",X"50",X"AB",X"80",X"97",X"50",X"39",X"D6",X"4F",
		X"EB",X"80",X"D7",X"51",X"39",X"D6",X"51",X"EB",X"80",X"D7",X"51",X"39",X"EC",X"81",X"DD",X"4E",
		X"DD",X"50",X"39",X"96",X"4E",X"D6",X"51",X"DB",X"4D",X"DD",X"50",X"39",X"10",X"AE",X"81",X"9F",
		X"52",X"9E",X"3D",X"AD",X"84",X"AB",X"A4",X"9B",X"4C",X"97",X"50",X"32",X"62",X"9E",X"3F",X"6E",
		X"84",X"34",X"77",X"10",X"8E",X"FF",X"B3",X"CE",X"CC",X"0F",X"20",X"1F",X"34",X"77",X"10",X"8E",
		X"FF",X"B6",X"CE",X"CC",X"0F",X"20",X"14",X"34",X"77",X"10",X"8E",X"FF",X"B3",X"CE",X"CC",X"39",
		X"20",X"09",X"34",X"77",X"10",X"8E",X"FF",X"B6",X"CE",X"CC",X"39",X"10",X"9F",X"3D",X"DF",X"3F",
		X"DE",X"59",X"11",X"83",X"FF",X"FF",X"26",X"15",X"9F",X"50",X"DD",X"59",X"26",X"05",X"CC",X"0F",
		X"FF",X"20",X"08",X"85",X"F0",X"26",X"04",X"8D",X"35",X"20",X"F8",X"DD",X"59",X"DC",X"59",X"84",
		X"F0",X"81",X"F0",X"26",X"07",X"35",X"77",X"9E",X"50",X"1A",X"01",X"39",X"44",X"44",X"8E",X"C5",
		X"FB",X"31",X"86",X"DC",X"50",X"9E",X"3D",X"AD",X"84",X"AB",X"A4",X"9B",X"4C",X"97",X"50",X"DC",
		X"59",X"8D",X"0B",X"DD",X"59",X"9E",X"3F",X"6E",X"84",X"35",X"77",X"1C",X"FE",X"39",X"58",X"49",
		X"58",X"49",X"58",X"49",X"58",X"49",X"CA",X"0F",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"38",X"4E",X"CE",X"96",X"09",X"AC",X"42",X"90",X"16",X"52",X"A8",X"F2",X"12",X"96",X"6A",
		X"08",X"C0",X"DE",X"CA",X"A5",X"54",X"1B",X"88",X"2D",X"59",X"A3",X"96",X"41",X"DC",X"EF",X"A3",
		X"27",X"03",X"B6",X"1C",X"EF",X"5E",X"FF",X"D7",X"B0",X"56",X"A4",X"76",X"C3",X"A0",X"90",X"9B",
		X"D9",X"08",X"D3",X"04",X"CB",X"99",X"C8",X"70",X"43",X"94",X"33",X"7B",X"6B",X"8D",X"B2",X"F8",
		X"00",X"0C",X"CC",X"CC",X"CC",X"CC",X"0C",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"C0",X"CC",X"CC",X"CC",X"CC",X"C0",X"00",
		X"A0",X"0A",X"A0",X"A0",X"00",X"A0",X"0A",X"00",X"0A",X"0A",X"A0",X"0A",X"0A",X"AA",X"0A",X"00",
		X"A0",X"00",X"00",X"0A",X"00",X"A0",X"AA",X"A0",X"00",X"02",X"23",X"02",X"20",X"22",X"23",X"22",
		X"00",X"00",X"20",X"00",X"00",X"00",X"02",X"00",X"02",X"22",X"32",X"22",X"00",X"20",X"32",X"20",
		X"00",X"00",X"03",X"03",X"00",X"00",X"03",X"30",X"04",X"34",X"30",X"30",X"34",X"30",X"00",X"00",
		X"44",X"44",X"33",X"33",X"34",X"30",X"30",X"30",X"00",X"30",X"03",X"03",X"30",X"30",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"03",X"33",X"33",X"03",X"03",X"30",X"00",X"44",X"44",X"03",X"03",X"43",X"03",X"03",X"03",
		X"40",X"43",X"30",X"30",X"43",X"03",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"30",X"03",
		X"00",X"00",X"03",X"03",X"00",X"00",X"03",X"30",X"04",X"34",X"03",X"03",X"34",X"30",X"00",X"00",
		X"44",X"44",X"30",X"30",X"34",X"30",X"30",X"30",X"00",X"30",X"33",X"33",X"30",X"30",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"03",X"30",X"30",X"03",X"03",X"30",X"00",X"44",X"44",X"33",X"33",X"43",X"03",X"03",X"03",
		X"40",X"43",X"03",X"03",X"43",X"03",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"30",X"03",
		X"00",X"00",X"03",X"03",X"00",X"00",X"03",X"30",X"00",X"33",X"33",X"33",X"33",X"30",X"00",X"00",
		X"00",X"33",X"03",X"03",X"33",X"30",X"30",X"30",X"00",X"30",X"33",X"33",X"30",X"30",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"03",X"33",X"33",X"03",X"03",X"30",X"00",X"00",X"33",X"30",X"30",X"03",X"03",X"03",X"03",
		X"00",X"33",X"33",X"33",X"33",X"03",X"00",X"00",X"00",X"00",X"30",X"30",X"00",X"00",X"30",X"03",
		X"00",X"03",X"34",X"03",X"33",X"70",X"40",X"33",X"33",X"07",X"44",X"33",X"33",X"00",X"04",X"33",
		X"30",X"73",X"40",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",X"00",X"03",X"37",X"44",X"33",
		X"33",X"00",X"04",X"33",X"33",X"70",X"40",X"33",X"33",X"07",X"44",X"33",X"00",X"30",X"03",X"30",
		X"00",X"03",X"30",X"03",X"33",X"00",X"44",X"33",X"33",X"70",X"04",X"33",X"33",X"07",X"40",X"33",
		X"30",X"03",X"44",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",X"00",X"03",X"30",X"04",X"33",
		X"33",X"07",X"40",X"33",X"33",X"00",X"44",X"33",X"33",X"70",X"04",X"33",X"00",X"30",X"43",X"30",
		X"00",X"03",X"34",X"03",X"33",X"07",X"04",X"33",X"33",X"00",X"40",X"33",X"33",X"70",X"44",X"33",
		X"30",X"03",X"04",X"33",X"00",X"00",X"30",X"00",X"00",X"00",X"03",X"00",X"03",X"30",X"40",X"33",
		X"33",X"70",X"44",X"33",X"33",X"07",X"04",X"33",X"33",X"00",X"40",X"33",X"00",X"30",X"43",X"30",
		X"00",X"06",X"26",X"06",X"26",X"00",X"66",X"66",X"66",X"88",X"88",X"88",X"00",X"60",X"66",X"66",
		X"88",X"86",X"00",X"00",X"00",X"66",X"66",X"93",X"00",X"00",X"00",X"6D",X"66",X"00",X"00",X"00",
		X"00",X"EF",X"66",X"00",X"00",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"02",X"00",X"02",X"00",X"06",X"66",X"66",X"28",X"68",X"08",X"60",X"66",X"66",X"86",
		X"88",X"88",X"00",X"00",X"60",X"66",X"86",X"69",X"00",X"00",X"00",X"66",X"66",X"30",X"00",X"00",
		X"00",X"DE",X"66",X"00",X"00",X"00",X"00",X"F0",X"66",X"00",X"00",X"00",X"00",X"00",X"93",X"00",
		X"00",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"00",X"0F",X"66",X"00",X"00",X"00",X"00",X"ED",
		X"66",X"00",X"00",X"00",X"00",X"66",X"66",X"03",X"00",X"00",X"06",X"66",X"68",X"96",X"06",X"66",
		X"66",X"68",X"88",X"88",X"60",X"66",X"66",X"83",X"86",X"80",X"00",X"00",X"30",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"00",X"FE",
		X"66",X"00",X"00",X"00",X"00",X"D6",X"66",X"00",X"00",X"00",X"00",X"66",X"66",X"39",X"00",X"06",
		X"66",X"66",X"88",X"68",X"66",X"66",X"66",X"88",X"88",X"88",X"00",X"60",X"63",X"30",X"63",X"00",
		X"06",X"26",X"68",X"28",X"60",X"66",X"66",X"86",X"00",X"00",X"66",X"66",X"00",X"00",X"ED",X"66",
		X"00",X"00",X"00",X"63",X"90",X"09",X"90",X"99",X"99",X"99",X"90",X"CC",X"90",X"11",X"00",X"11",
		X"10",X"11",X"00",X"10",X"10",X"10",X"00",X"10",X"00",X"11",X"10",X"11",X"00",X"11",X"00",X"10",
		X"00",X"10",X"10",X"10",X"00",X"11",X"10",X"10",X"10",X"11",X"00",X"10",X"10",X"10",X"10",X"10",
		X"00",X"01",X"00",X"01",X"01",X"01",X"00",X"11",X"01",X"11",X"00",X"11",X"00",X"01",X"01",X"01",
		X"00",X"01",X"00",X"11",X"00",X"11",X"01",X"11",X"00",X"01",X"01",X"01",X"01",X"01",X"00",X"11",
		X"01",X"01",X"01",X"11",X"00",X"FF",X"F0",X"FF",X"00",X"FF",X"00",X"F0",X"00",X"F0",X"F0",X"F0",
		X"00",X"EE",X"E0",X"E0",X"E0",X"EE",X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"DD",X"D0",X"D0",
		X"D0",X"DD",X"00",X"D0",X"D0",X"D0",X"D0",X"D0",X"00",X"0F",X"0F",X"0F",X"00",X"0F",X"00",X"FF",
		X"00",X"FF",X"0F",X"FF",X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"EE",X"0E",X"0E",X"0E",X"EE",
		X"00",X"0D",X"0D",X"0D",X"0D",X"0D",X"00",X"DD",X"0D",X"0D",X"0D",X"DD",X"00",X"1C",X"0D",X"7F",
		X"E7",X"70",X"00",X"0F",X"71",X"71",X"07",X"DC",X"77",X"7C",X"0D",X"71",X"C7",X"77",X"DE",X"07",
		X"71",X"17",X"17",X"DE",X"F7",X"71",X"17",X"71",X"7C",X"DE",X"F0",X"07",X"77",X"C7",X"71",X"17",
		X"70",X"70",X"7C",X"D7",X"77",X"77",X"70",X"01",X"CD",X"FF",X"D7",X"70",X"F0",X"00",X"00",X"00",
		X"7E",X"C0",X"76",X"7E",X"C0",X"9C",X"7E",X"C0",X"B8",X"7E",X"C0",X"FC",X"7E",X"CB",X"E6",X"7E",
		X"CB",X"E0",X"7E",X"CC",X"2C",X"7E",X"CC",X"20",X"7E",X"CC",X"26",X"7E",X"CC",X"AF",X"7E",X"CB",
		X"AF",X"7E",X"C7",X"99",X"7E",X"C1",X"27",X"7E",X"C1",X"46",X"7E",X"C2",X"3D",X"7E",X"C2",X"C3",
		X"7E",X"C4",X"06",X"7E",X"CC",X"C1",X"7E",X"FF",X"D4",X"7E",X"FF",X"D7",X"BD",X"FF",X"CE",X"C0",
		X"02",X"02",X"39",X"BD",X"FF",X"CE",X"C0",X"05",X"02",X"39",X"BD",X"FF",X"CE",X"C0",X"0E",X"02",
		X"39",X"BD",X"FF",X"CE",X"C0",X"11",X"02",X"39",X"BD",X"FF",X"CE",X"C0",X"1A",X"02",X"39",X"BD",
		X"FF",X"CE",X"C0",X"1D",X"02",X"39",X"BD",X"FF",X"CE",X"C0",X"20",X"02",X"39",X"BD",X"FF",X"CE",
		X"C0",X"23",X"02",X"39",X"D9",X"FF",X"BD",X"CA",X"2A",X"C6",X"7A",X"BD",X"C7",X"93",X"CE",X"C0",
		X"69",X"8E",X"28",X"70",X"BD",X"C0",X"3C",X"CE",X"C0",X"6B",X"8E",X"40",X"90",X"BD",X"C0",X"3C",
		X"C6",X"0F",X"BD",X"CA",X"C8",X"10",X"8E",X"0B",X"B8",X"7E",X"CA",X"44",X"BD",X"CA",X"2A",X"C6",
		X"57",X"BD",X"C7",X"93",X"CE",X"C0",X"69",X"8E",X"28",X"70",X"BD",X"C0",X"3C",X"CE",X"C0",X"73",
		X"8E",X"38",X"90",X"BD",X"C0",X"3C",X"20",X"29",X"BD",X"CA",X"2A",X"C6",X"57",X"BD",X"C7",X"93",
		X"CE",X"C0",X"69",X"8E",X"28",X"60",X"BD",X"C0",X"3C",X"CE",X"C0",X"71",X"8E",X"38",X"80",X"BD",
		X"C0",X"3C",X"1F",X"B8",X"81",X"9E",X"27",X"09",X"CE",X"C0",X"73",X"8E",X"38",X"A0",X"BD",X"C0",
		X"3C",X"10",X"8E",X"0B",X"B8",X"BD",X"CA",X"57",X"8E",X"CC",X"00",X"BD",X"C0",X"39",X"C5",X"02",
		X"27",X"05",X"54",X"25",X"06",X"20",X"4F",X"31",X"3F",X"26",X"EA",X"39",X"1C",X"EF",X"8E",X"C4",
		X"7F",X"BD",X"FF",X"A4",X"C1",X"5A",X"26",X"36",X"8E",X"C4",X"00",X"BD",X"C0",X"39",X"C4",X"0F",
		X"26",X"01",X"39",X"5F",X"BD",X"C0",X"36",X"8E",X"C4",X"7D",X"BD",X"FF",X"A4",X"4F",X"30",X"1E",
		X"BD",X"FF",X"AA",X"C1",X"15",X"26",X"04",X"1C",X"7F",X"20",X"1B",X"C1",X"25",X"26",X"03",X"7E",
		X"CC",X"AF",X"C1",X"35",X"26",X"03",X"7E",X"CB",X"BF",X"C1",X"45",X"27",X"01",X"39",X"32",X"62",
		X"BD",X"CB",X"CF",X"7E",X"C7",X"99",X"1A",X"10",X"BD",X"CA",X"2A",X"BD",X"FF",X"BF",X"34",X"40",
		X"FE",X"FF",X"9F",X"33",X"C8",X"18",X"DF",X"43",X"35",X"40",X"11",X"93",X"43",X"27",X"70",X"DF",
		X"5B",X"C6",X"08",X"BD",X"CA",X"AA",X"C6",X"57",X"BD",X"C7",X"93",X"CE",X"C0",X"71",X"8E",X"38",
		X"60",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",X"35",X"BD",X"C0",X"6D",X"CC",X"42",X"66",X"DD",X"4A",
		X"9E",X"4A",X"30",X"0A",X"9F",X"4A",X"CE",X"C0",X"6D",X"BD",X"C0",X"3C",X"FE",X"FF",X"9F",X"DF",
		X"43",X"DE",X"5B",X"DC",X"5B",X"93",X"43",X"54",X"25",X"02",X"33",X"41",X"5C",X"D7",X"3A",X"BD",
		X"CB",X"23",X"9E",X"50",X"BD",X"C0",X"4A",X"BD",X"CA",X"69",X"BD",X"FF",X"C2",X"DF",X"5B",X"FE",
		X"FF",X"9F",X"33",X"C8",X"18",X"11",X"93",X"5B",X"26",X"C6",X"BD",X"CA",X"0E",X"0D",X"49",X"26",
		X"30",X"D6",X"3A",X"BD",X"CA",X"AA",X"10",X"8E",X"C0",X"39",X"BD",X"C0",X"6D",X"20",X"1F",X"1F",
		X"A9",X"5D",X"2A",X"3E",X"C6",X"7A",X"BD",X"C7",X"93",X"CE",X"C0",X"77",X"8E",X"38",X"80",X"BD",
		X"C0",X"3C",X"10",X"8E",X"C0",X"39",X"BD",X"C0",X"6D",X"C6",X"08",X"BD",X"CA",X"C8",X"BD",X"CA",
		X"39",X"BD",X"CA",X"2A",X"5F",X"BD",X"CA",X"AA",X"BD",X"C7",X"91",X"CE",X"C0",X"79",X"8E",X"40",
		X"80",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",X"3D",X"BD",X"C0",X"6D",X"10",X"8E",X"13",X"88",X"BD",
		X"CA",X"44",X"BD",X"CA",X"57",X"0D",X"49",X"10",X"26",X"00",X"D7",X"0D",X"47",X"26",X"F3",X"8E",
		X"C0",X"00",X"C6",X"C0",X"BD",X"C0",X"36",X"86",X"B5",X"3D",X"1E",X"89",X"30",X"01",X"8C",X"C0",
		X"10",X"26",X"F1",X"CC",X"00",X"00",X"10",X"8E",X"00",X"0A",X"7E",X"FF",X"C5",X"1F",X"20",X"E8",
		X"82",X"A8",X"82",X"DD",X"41",X"9F",X"43",X"BD",X"CA",X"F9",X"BD",X"FF",X"BC",X"BD",X"CA",X"E4",
		X"BD",X"CA",X"69",X"C6",X"04",X"BD",X"CA",X"AA",X"C6",X"57",X"BD",X"C7",X"93",X"CE",X"C0",X"73",
		X"8E",X"38",X"70",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",X"41",X"BD",X"C0",X"6D",X"DC",X"41",X"4D",
		X"26",X"02",X"1F",X"98",X"5F",X"5C",X"44",X"24",X"FC",X"D7",X"3A",X"DC",X"43",X"80",X"03",X"24",
		X"FC",X"8B",X"04",X"97",X"3B",X"CE",X"C0",X"6F",X"8E",X"42",X"90",X"BD",X"C0",X"3C",X"D6",X"3B",
		X"58",X"58",X"58",X"58",X"DB",X"3A",X"4F",X"9E",X"50",X"BD",X"C0",X"4A",X"BD",X"CA",X"0E",X"0D",
		X"49",X"26",X"4F",X"96",X"3B",X"C6",X"10",X"54",X"4A",X"26",X"FC",X"BD",X"CA",X"AA",X"BD",X"CA",
		X"0E",X"0D",X"49",X"26",X"3D",X"D6",X"3A",X"BD",X"CA",X"AA",X"10",X"8E",X"C0",X"45",X"BD",X"C0",
		X"6D",X"20",X"2C",X"BD",X"CA",X"F9",X"BD",X"FF",X"BC",X"BD",X"CA",X"E4",X"BD",X"CA",X"69",X"10",
		X"8C",X"00",X"0A",X"27",X"1D",X"C6",X"7A",X"BD",X"C7",X"93",X"CE",X"C0",X"7B",X"8E",X"28",X"80",
		X"BD",X"C0",X"3C",X"10",X"8E",X"C0",X"45",X"BD",X"C0",X"6D",X"C6",X"04",X"BD",X"CA",X"C8",X"BD",
		X"CA",X"39",X"BD",X"CA",X"2A",X"1F",X"B8",X"81",X"A2",X"26",X"1D",X"C6",X"02",X"BD",X"CA",X"AA",
		X"C6",X"57",X"BD",X"C7",X"93",X"CE",X"C0",X"81",X"8E",X"28",X"80",X"BD",X"C0",X"3C",X"10",X"8E",
		X"C0",X"49",X"BD",X"C0",X"6D",X"7E",X"C3",X"BB",X"8B",X"03",X"5F",X"DD",X"41",X"DE",X"41",X"8E",
		X"C4",X"00",X"BD",X"C0",X"39",X"E7",X"C0",X"30",X"01",X"8C",X"C5",X"00",X"26",X"F4",X"CC",X"00",
		X"10",X"D7",X"3A",X"4F",X"8E",X"C4",X"00",X"D6",X"3A",X"BD",X"C0",X"36",X"30",X"01",X"5C",X"D1",
		X"3A",X"26",X"F6",X"8E",X"C4",X"00",X"4C",X"BD",X"C0",X"39",X"D7",X"3B",X"30",X"01",X"BD",X"C0",
		X"39",X"D0",X"3B",X"5A",X"C4",X"0F",X"26",X"0E",X"4C",X"26",X"EC",X"BD",X"CA",X"69",X"0D",X"49",
		X"26",X"04",X"0A",X"3A",X"26",X"CE",X"DE",X"41",X"8E",X"C4",X"00",X"E6",X"C0",X"BD",X"C0",X"36",
		X"30",X"01",X"8C",X"C5",X"00",X"26",X"F4",X"0D",X"49",X"26",X"43",X"96",X"3A",X"27",X"22",X"C6",
		X"02",X"BD",X"CA",X"AA",X"C6",X"57",X"BD",X"C7",X"93",X"BD",X"CA",X"69",X"CE",X"C0",X"7D",X"8E",
		X"30",X"80",X"BD",X"C0",X"3C",X"BD",X"CA",X"69",X"10",X"8E",X"C0",X"49",X"BD",X"C0",X"6D",X"20",
		X"1A",X"C6",X"7A",X"BD",X"C7",X"93",X"CE",X"C0",X"7F",X"8E",X"38",X"80",X"BD",X"C0",X"3C",X"10",
		X"8E",X"C0",X"49",X"BD",X"C0",X"6D",X"C6",X"02",X"BD",X"CA",X"C8",X"BD",X"CA",X"39",X"BD",X"CA",
		X"2A",X"C6",X"01",X"BD",X"CA",X"AA",X"BD",X"C7",X"91",X"CE",X"C0",X"83",X"8E",X"38",X"80",X"BD",
		X"C0",X"3C",X"10",X"8E",X"C0",X"4D",X"BD",X"C0",X"6D",X"10",X"8E",X"13",X"88",X"BD",X"CA",X"44",
		X"BD",X"CB",X"67",X"10",X"8E",X"07",X"D0",X"CE",X"C9",X"D8",X"E6",X"C0",X"8E",X"C0",X"00",X"BD",
		X"C0",X"36",X"30",X"01",X"8C",X"C0",X"10",X"26",X"F6",X"BD",X"CA",X"44",X"11",X"83",X"C9",X"E0",
		X"26",X"E8",X"0D",X"49",X"27",X"E1",X"BD",X"CA",X"2A",X"5F",X"D7",X"41",X"D7",X"42",X"BD",X"CA",
		X"AA",X"BD",X"C7",X"91",X"CE",X"C0",X"85",X"8E",X"40",X"78",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",
		X"55",X"BD",X"C0",X"6D",X"10",X"8E",X"00",X"01",X"CE",X"C9",X"F0",X"4F",X"8E",X"CC",X"00",X"BD",
		X"C0",X"39",X"C5",X"01",X"26",X"09",X"C5",X"02",X"26",X"15",X"BD",X"CA",X"57",X"20",X"ED",X"BD",
		X"CA",X"44",X"4C",X"A1",X"C4",X"26",X"04",X"33",X"41",X"20",X"F7",X"97",X"3A",X"88",X"3F",X"C6",
		X"13",X"BD",X"CB",X"0B",X"0D",X"49",X"26",X"2E",X"D6",X"3A",X"BD",X"CB",X"0B",X"10",X"8E",X"03",
		X"E8",X"DC",X"41",X"8E",X"5A",X"8C",X"BD",X"C0",X"51",X"D6",X"3A",X"BD",X"CB",X"23",X"4F",X"DD",
		X"41",X"8E",X"5A",X"8C",X"BD",X"C0",X"4A",X"96",X"3A",X"81",X"1F",X"26",X"AF",X"1F",X"A9",X"5D",
		X"10",X"2A",X"01",X"01",X"20",X"A2",X"BD",X"CA",X"2A",X"BD",X"C7",X"91",X"CE",X"C0",X"87",X"8E",
		X"38",X"20",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",X"59",X"BD",X"C0",X"6D",X"1F",X"B8",X"C6",X"62",
		X"DD",X"41",X"CB",X"26",X"1F",X"01",X"86",X"FF",X"A7",X"82",X"9C",X"41",X"26",X"FA",X"0F",X"5D",
		X"0F",X"5E",X"0F",X"5F",X"0F",X"60",X"0F",X"61",X"86",X"01",X"97",X"3C",X"8E",X"CC",X"00",X"DE",
		X"41",X"33",X"5B",X"4F",X"BD",X"C0",X"39",X"8C",X"CC",X"06",X"26",X"02",X"C4",X"7F",X"81",X"18",
		X"26",X"02",X"C4",X"CF",X"D7",X"3A",X"E8",X"C0",X"26",X"38",X"8B",X"08",X"30",X"02",X"8C",X"CC",
		X"02",X"27",X"F9",X"8C",X"CC",X"08",X"26",X"DC",X"81",X"28",X"27",X"15",X"30",X"1E",X"BD",X"C0",
		X"39",X"5D",X"2A",X"0D",X"C6",X"34",X"30",X"01",X"BD",X"C0",X"36",X"30",X"1D",X"0C",X"3C",X"20",
		X"C3",X"C6",X"3C",X"8E",X"CC",X"07",X"BD",X"C0",X"36",X"BD",X"CA",X"69",X"0D",X"49",X"27",X"A8",
		X"20",X"73",X"D7",X"3B",X"C6",X"01",X"D5",X"3B",X"26",X"04",X"4C",X"58",X"20",X"F8",X"9E",X"41",
		X"D5",X"3A",X"26",X"14",X"E8",X"C2",X"E7",X"C4",X"A1",X"80",X"26",X"FC",X"63",X"82",X"8D",X"3C",
		X"CC",X"38",X"08",X"BD",X"FF",X"B9",X"20",X"C9",X"E8",X"C2",X"E7",X"C4",X"C6",X"08",X"BD",X"CB",
		X"0B",X"6D",X"80",X"2A",X"FC",X"A7",X"82",X"34",X"02",X"8D",X"21",X"BD",X"C0",X"3C",X"35",X"02",
		X"81",X"08",X"25",X"AD",X"44",X"81",X"06",X"27",X"A8",X"8E",X"CC",X"06",X"BD",X"C0",X"39",X"5D",
		X"2A",X"9F",X"9E",X"50",X"4F",X"D6",X"3C",X"BD",X"C0",X"4A",X"20",X"95",X"CE",X"C0",X"8B",X"81",
		X"18",X"25",X"02",X"80",X"10",X"48",X"33",X"C6",X"1F",X"10",X"93",X"41",X"86",X"0A",X"3D",X"C3",
		X"38",X"30",X"1F",X"01",X"39",X"BD",X"CA",X"2A",X"BD",X"C7",X"91",X"CE",X"C0",X"89",X"8E",X"28",
		X"80",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",X"5D",X"BD",X"C0",X"6D",X"8E",X"CC",X"00",X"CE",X"C9",
		X"F4",X"BD",X"C0",X"39",X"C5",X"01",X"27",X"14",X"10",X"8E",X"13",X"88",X"BD",X"CA",X"44",X"0D",
		X"49",X"10",X"26",X"01",X"E4",X"BD",X"C0",X"39",X"C5",X"01",X"26",X"09",X"BD",X"CA",X"0E",X"0D",
		X"49",X"10",X"26",X"01",X"D4",X"34",X"70",X"AD",X"D4",X"35",X"70",X"33",X"42",X"11",X"83",X"C9",
		X"FE",X"26",X"CE",X"10",X"8E",X"13",X"88",X"BD",X"CA",X"44",X"1F",X"A9",X"5D",X"10",X"2A",X"FB",
		X"65",X"20",X"BB",X"BD",X"CA",X"69",X"BD",X"FF",X"BC",X"BD",X"CA",X"F9",X"8E",X"C0",X"01",X"C6",
		X"FF",X"BD",X"C0",X"36",X"8E",X"C0",X"02",X"C6",X"C0",X"BD",X"C0",X"36",X"8E",X"C0",X"03",X"C6",
		X"38",X"BD",X"C0",X"36",X"8E",X"C0",X"04",X"C6",X"07",X"BD",X"C0",X"36",X"BD",X"CA",X"69",X"10",
		X"8E",X"C6",X"F7",X"CC",X"01",X"01",X"AE",X"A4",X"ED",X"81",X"AC",X"22",X"26",X"FA",X"31",X"24",
		X"10",X"8C",X"C7",X"1F",X"26",X"F0",X"BD",X"CA",X"69",X"86",X"11",X"10",X"8E",X"C6",X"D7",X"AE",
		X"A4",X"9F",X"45",X"A7",X"84",X"0C",X"45",X"9E",X"45",X"AC",X"22",X"26",X"F6",X"31",X"24",X"10",
		X"8C",X"C6",X"F7",X"26",X"EA",X"BD",X"CA",X"69",X"10",X"8E",X"C7",X"1F",X"AE",X"A4",X"9F",X"45",
		X"A6",X"24",X"A7",X"84",X"0C",X"45",X"9E",X"45",X"AC",X"22",X"26",X"F6",X"31",X"25",X"10",X"8C",
		X"C7",X"5B",X"26",X"E8",X"BD",X"CA",X"69",X"10",X"8E",X"C7",X"5B",X"AE",X"A4",X"A6",X"24",X"A7",
		X"80",X"AC",X"22",X"26",X"FA",X"31",X"25",X"10",X"8C",X"C7",X"6F",X"26",X"EE",X"BD",X"CA",X"69",
		X"86",X"21",X"B7",X"46",X"7E",X"86",X"20",X"B7",X"96",X"7E",X"8E",X"4E",X"0A",X"A6",X"84",X"84",
		X"F0",X"8A",X"02",X"A7",X"80",X"8C",X"4E",X"6D",X"26",X"F3",X"8E",X"4E",X"90",X"A6",X"84",X"84",
		X"F0",X"8A",X"02",X"A7",X"80",X"8C",X"4E",X"F3",X"26",X"F3",X"BD",X"CA",X"69",X"8E",X"0E",X"18",
		X"9F",X"45",X"9E",X"45",X"A6",X"84",X"84",X"F0",X"8A",X"01",X"A7",X"84",X"D6",X"46",X"CB",X"22",
		X"25",X"04",X"D7",X"46",X"20",X"EC",X"C6",X"18",X"D7",X"46",X"D6",X"45",X"CB",X"10",X"D7",X"45",
		X"C1",X"9E",X"26",X"DE",X"7E",X"CA",X"69",X"07",X"07",X"97",X"07",X"07",X"29",X"97",X"29",X"07",
		X"4B",X"97",X"4B",X"07",X"6D",X"97",X"6D",X"07",X"8F",X"97",X"8F",X"07",X"B1",X"97",X"B1",X"07",
		X"D3",X"97",X"D3",X"07",X"F5",X"97",X"F5",X"06",X"07",X"06",X"F5",X"16",X"07",X"16",X"F5",X"26",
		X"07",X"26",X"F5",X"36",X"07",X"36",X"F5",X"46",X"07",X"46",X"F5",X"56",X"07",X"56",X"F5",X"66",
		X"07",X"66",X"F5",X"76",X"07",X"76",X"F5",X"86",X"07",X"86",X"F5",X"96",X"07",X"96",X"F5",X"48",
		X"05",X"55",X"05",X"44",X"48",X"06",X"55",X"06",X"44",X"48",X"07",X"55",X"07",X"00",X"48",X"08",
		X"55",X"08",X"33",X"48",X"09",X"55",X"09",X"33",X"48",X"F3",X"55",X"F3",X"33",X"48",X"F4",X"55",
		X"F4",X"33",X"48",X"F5",X"55",X"F5",X"00",X"48",X"F6",X"55",X"F6",X"44",X"48",X"F7",X"55",X"F7",
		X"44",X"07",X"7E",X"46",X"7E",X"22",X"57",X"7E",X"96",X"7E",X"22",X"05",X"6F",X"05",X"8E",X"04",
		X"06",X"6F",X"06",X"8E",X"30",X"96",X"6F",X"96",X"8E",X"00",X"97",X"6F",X"97",X"8E",X"34",X"BD",
		X"FF",X"BC",X"C6",X"05",X"8E",X"C0",X"00",X"8D",X"03",X"8E",X"C0",X"0C",X"7E",X"C0",X"36",X"C6",
		X"28",X"20",X"F1",X"C6",X"80",X"20",X"ED",X"10",X"8E",X"C9",X"FE",X"BD",X"CA",X"97",X"7E",X"CB",
		X"3B",X"C6",X"A5",X"8E",X"C0",X"01",X"7E",X"C0",X"36",X"BD",X"CA",X"69",X"BD",X"CA",X"2A",X"8D",
		X"F0",X"CE",X"C0",X"D7",X"8E",X"28",X"20",X"BD",X"CA",X"69",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",
		X"61",X"BD",X"C0",X"6D",X"10",X"8E",X"05",X"DC",X"BD",X"CA",X"44",X"0D",X"49",X"26",X"60",X"0F",
		X"3C",X"86",X"01",X"97",X"3B",X"32",X"E8",X"E0",X"BD",X"FF",X"BC",X"CE",X"C0",X"D7",X"8E",X"28",
		X"20",X"BD",X"CA",X"69",X"BD",X"C0",X"3C",X"0F",X"3A",X"10",X"8E",X"C0",X"65",X"BD",X"C0",X"66",
		X"BD",X"CA",X"69",X"86",X"20",X"1F",X"89",X"5A",X"30",X"E4",X"A7",X"80",X"5A",X"26",X"FB",X"86",
		X"2F",X"A7",X"80",X"30",X"E4",X"BD",X"CA",X"57",X"8E",X"CC",X"00",X"BD",X"C0",X"39",X"C5",X"02",
		X"27",X"23",X"C5",X"01",X"26",X"0C",X"0C",X"3B",X"0A",X"3C",X"2A",X"19",X"C6",X"1B",X"D7",X"3C",
		X"20",X"13",X"0C",X"3C",X"0C",X"3B",X"86",X"1C",X"91",X"3C",X"26",X"09",X"32",X"E8",X"20",X"BD",
		X"CA",X"69",X"7E",X"FF",X"C8",X"BD",X"C9",X"7A",X"0D",X"3B",X"27",X"C9",X"D6",X"3C",X"C1",X"09",
		X"26",X"25",X"8E",X"C4",X"87",X"BD",X"FF",X"A4",X"5D",X"27",X"1C",X"C1",X"08",X"22",X"05",X"BD",
		X"CB",X"99",X"20",X"13",X"8E",X"C4",X"87",X"34",X"10",X"C6",X"01",X"BD",X"FF",X"AD",X"BD",X"CB",
		X"99",X"5F",X"35",X"10",X"BD",X"FF",X"AD",X"8D",X"38",X"96",X"3A",X"81",X"06",X"27",X"0E",X"4D",
		X"26",X"04",X"86",X"64",X"20",X"02",X"86",X"06",X"97",X"3A",X"4C",X"C6",X"FF",X"BD",X"CA",X"57",
		X"4A",X"27",X"19",X"8E",X"CC",X"00",X"34",X"04",X"BD",X"C0",X"39",X"C5",X"0A",X"26",X"04",X"1C",
		X"FE",X"20",X"02",X"1A",X"01",X"35",X"04",X"56",X"26",X"E3",X"0F",X"3A",X"0F",X"3B",X"7E",X"C7",
		X"F5",X"31",X"62",X"8E",X"10",X"80",X"BD",X"C0",X"58",X"BD",X"C9",X"1F",X"96",X"3C",X"4C",X"BD",
		X"C9",X"02",X"BD",X"C9",X"10",X"ED",X"84",X"D6",X"3C",X"58",X"58",X"8E",X"CC",X"D6",X"3A",X"10",
		X"AE",X"84",X"EE",X"02",X"30",X"6E",X"A6",X"A0",X"81",X"2F",X"27",X"04",X"A7",X"80",X"20",X"F6",
		X"1F",X"30",X"33",X"62",X"8E",X"C4",X"00",X"3A",X"BD",X"FF",X"A4",X"34",X"06",X"D6",X"3C",X"5C",
		X"C1",X"07",X"22",X"13",X"35",X"06",X"1F",X"98",X"BD",X"C9",X"10",X"ED",X"47",X"BD",X"FF",X"A1",
		X"BD",X"C9",X"10",X"ED",X"49",X"20",X"13",X"C1",X"08",X"26",X"09",X"CC",X"30",X"30",X"ED",X"49",
		X"33",X"5E",X"20",X"E0",X"35",X"06",X"1F",X"98",X"20",X"E6",X"8E",X"10",X"80",X"31",X"62",X"7E",
		X"C0",X"5F",X"34",X"04",X"1F",X"89",X"86",X"99",X"8B",X"01",X"19",X"5A",X"2A",X"FA",X"35",X"84",
		X"1F",X"89",X"84",X"F0",X"44",X"44",X"44",X"44",X"8B",X"30",X"C4",X"0F",X"CB",X"30",X"39",X"86",
		X"20",X"1F",X"89",X"5A",X"30",X"64",X"A7",X"80",X"5A",X"26",X"FB",X"86",X"2F",X"A7",X"80",X"30",
		X"64",X"39",X"8C",X"C4",X"81",X"26",X"1A",X"BD",X"FF",X"A7",X"30",X"1C",X"1E",X"89",X"8B",X"10",
		X"19",X"24",X"07",X"1E",X"89",X"8B",X"01",X"19",X"1E",X"89",X"1E",X"89",X"0C",X"3B",X"7E",X"FF",
		X"B0",X"BD",X"FF",X"A1",X"8B",X"01",X"19",X"30",X"1E",X"0C",X"3B",X"7E",X"FF",X"AA",X"8C",X"C4",
		X"81",X"26",X"10",X"BD",X"FF",X"A7",X"30",X"1C",X"1E",X"89",X"8B",X"90",X"19",X"1E",X"89",X"89",
		X"99",X"20",X"D4",X"BD",X"FF",X"A1",X"8B",X"99",X"20",X"DC",X"D6",X"3C",X"5C",X"C1",X"07",X"22",
		X"01",X"39",X"C1",X"09",X"23",X"11",X"C1",X"10",X"22",X"0D",X"C1",X"0A",X"27",X"09",X"8E",X"C4",
		X"87",X"BD",X"FF",X"A1",X"4D",X"26",X"EA",X"5A",X"58",X"58",X"8E",X"CC",X"D6",X"3A",X"E6",X"03",
		X"8E",X"C4",X"00",X"3A",X"34",X"10",X"BD",X"CA",X"57",X"8E",X"CC",X"00",X"BD",X"C0",X"39",X"C5",
		X"02",X"27",X"02",X"35",X"90",X"C5",X"08",X"26",X"04",X"0F",X"3A",X"20",X"E9",X"35",X"10",X"8C",
		X"C4",X"7D",X"26",X"0C",X"34",X"14",X"8E",X"C4",X"00",X"C6",X"01",X"BD",X"C0",X"36",X"35",X"14",
		X"54",X"10",X"25",X"FF",X"5D",X"7E",X"C9",X"5E",X"02",X"03",X"04",X"10",X"18",X"20",X"40",X"80",
		X"00",X"FF",X"11",X"EE",X"22",X"DD",X"33",X"CC",X"44",X"BB",X"55",X"AA",X"66",X"99",X"77",X"88",
		X"13",X"1B",X"1C",X"00",X"C5",X"E3",X"C7",X"6F",X"C7",X"7F",X"C7",X"83",X"C7",X"87",X"05",X"05",
		X"28",X"28",X"80",X"80",X"00",X"00",X"AD",X"AD",X"2D",X"2D",X"A8",X"A8",X"85",X"85",X"8E",X"CC",
		X"00",X"10",X"8E",X"00",X"64",X"BD",X"CA",X"44",X"BD",X"C0",X"39",X"C5",X"02",X"26",X"F6",X"BD",
		X"CA",X"44",X"BD",X"C0",X"39",X"C5",X"02",X"27",X"F6",X"39",X"BD",X"FF",X"BC",X"8D",X"3A",X"BD",
		X"CA",X"F9",X"0A",X"49",X"2A",X"02",X"0F",X"49",X"39",X"10",X"8E",X"00",X"01",X"8D",X"05",X"0D",
		X"49",X"27",X"FA",X"39",X"34",X"23",X"8D",X"21",X"0D",X"49",X"26",X"09",X"86",X"B2",X"4A",X"26",
		X"FD",X"31",X"3F",X"26",X"F1",X"35",X"A3",X"34",X"24",X"D6",X"49",X"0F",X"49",X"10",X"8E",X"00",
		X"0A",X"8D",X"E1",X"DB",X"49",X"D7",X"49",X"35",X"A4",X"34",X"15",X"C6",X"38",X"8E",X"C3",X"FC",
		X"BD",X"C0",X"36",X"8E",X"CC",X"00",X"BD",X"C0",X"39",X"53",X"C4",X"03",X"27",X"02",X"1C",X"FE",
		X"D6",X"47",X"56",X"D7",X"47",X"26",X"02",X"D7",X"48",X"53",X"26",X"09",X"D6",X"48",X"26",X"05",
		X"53",X"D7",X"48",X"0C",X"49",X"35",X"95",X"34",X"34",X"8E",X"C0",X"00",X"E6",X"A0",X"BD",X"C0",
		X"36",X"30",X"01",X"8C",X"C0",X"10",X"26",X"F4",X"35",X"B4",X"34",X"14",X"54",X"56",X"56",X"56",
		X"2A",X"01",X"5C",X"56",X"56",X"8E",X"CC",X"00",X"BD",X"C0",X"36",X"58",X"58",X"58",X"CA",X"3F",
		X"8E",X"CC",X"02",X"BD",X"C0",X"36",X"35",X"94",X"34",X"26",X"86",X"02",X"10",X"8E",X"01",X"F4",
		X"BD",X"CA",X"AA",X"BD",X"CA",X"44",X"5F",X"BD",X"CA",X"AA",X"BD",X"CA",X"44",X"E6",X"61",X"4A",
		X"26",X"EE",X"35",X"26",X"34",X"06",X"0F",X"52",X"0F",X"49",X"86",X"01",X"97",X"48",X"86",X"03",
		X"97",X"36",X"CC",X"FF",X"FF",X"DD",X"59",X"35",X"86",X"34",X"14",X"5F",X"8E",X"C0",X"00",X"BD",
		X"C0",X"36",X"30",X"01",X"8C",X"C0",X"10",X"26",X"F6",X"35",X"94",X"34",X"14",X"53",X"C4",X"3F",
		X"8E",X"CC",X"02",X"BD",X"C0",X"36",X"BD",X"CA",X"57",X"C6",X"3F",X"BD",X"C0",X"36",X"BD",X"CA",
		X"57",X"35",X"94",X"34",X"02",X"1F",X"98",X"84",X"0F",X"8B",X"00",X"19",X"C4",X"F0",X"27",X"07",
		X"8B",X"16",X"19",X"C0",X"10",X"20",X"F7",X"1F",X"89",X"35",X"82",X"34",X"16",X"CC",X"00",X"00",
		X"8E",X"00",X"00",X"9F",X"3D",X"30",X"89",X"0F",X"00",X"ED",X"83",X"9C",X"3D",X"26",X"FA",X"30",
		X"89",X"09",X"00",X"4D",X"26",X"03",X"8E",X"0F",X"00",X"BD",X"CA",X"69",X"0D",X"49",X"26",X"05",
		X"C3",X"11",X"11",X"24",X"DE",X"35",X"96",X"BD",X"CA",X"F9",X"8E",X"00",X"00",X"10",X"8E",X"C9",
		X"E0",X"9F",X"3D",X"30",X"89",X"0F",X"00",X"A6",X"A0",X"1F",X"89",X"ED",X"83",X"9C",X"3D",X"26",
		X"FA",X"30",X"89",X"09",X"00",X"4D",X"26",X"03",X"8E",X"0F",X"00",X"BD",X"CA",X"69",X"0D",X"49",
		X"26",X"06",X"10",X"8C",X"C9",X"F0",X"26",X"D9",X"39",X"8E",X"C4",X"87",X"BD",X"FF",X"AD",X"58",
		X"34",X"04",X"58",X"EB",X"E0",X"8E",X"CF",X"10",X"3A",X"10",X"8E",X"C4",X"89",X"C6",X"06",X"34",
		X"02",X"A6",X"80",X"1E",X"12",X"BD",X"FF",X"AA",X"1E",X"12",X"5A",X"26",X"F4",X"35",X"82",X"C6",
		X"0E",X"20",X"01",X"5F",X"8E",X"C4",X"00",X"4F",X"BD",X"FF",X"AA",X"5A",X"26",X"FA",X"39",X"34",
		X"36",X"8D",X"F0",X"8E",X"CE",X"CF",X"10",X"8E",X"C4",X"1D",X"C6",X"47",X"8D",X"D1",X"35",X"B6",
		X"34",X"16",X"86",X"01",X"20",X"02",X"34",X"16",X"C4",X"07",X"27",X"1F",X"58",X"58",X"8E",X"C3",
		X"FD",X"3A",X"BD",X"FF",X"A4",X"34",X"04",X"BD",X"FF",X"A4",X"34",X"04",X"AB",X"E0",X"19",X"1E",
		X"89",X"35",X"02",X"89",X"00",X"19",X"30",X"1C",X"BD",X"FF",X"B0",X"35",X"96",X"34",X"12",X"9B",
		X"37",X"19",X"24",X"02",X"86",X"99",X"97",X"37",X"8E",X"C4",X"7D",X"BD",X"FF",X"AA",X"35",X"92",
		X"34",X"16",X"C6",X"03",X"20",X"0A",X"34",X"16",X"C6",X"02",X"20",X"04",X"34",X"16",X"C6",X"01",
		X"BD",X"CB",X"E0",X"58",X"8E",X"C4",X"87",X"3A",X"BD",X"FF",X"A4",X"8D",X"62",X"96",X"39",X"34",
		X"04",X"AB",X"E4",X"97",X"39",X"96",X"38",X"AB",X"E0",X"97",X"38",X"8E",X"C4",X"93",X"BD",X"FF",
		X"A4",X"8D",X"4C",X"34",X"04",X"A1",X"E0",X"24",X"02",X"35",X"96",X"8E",X"C4",X"8F",X"BD",X"FF",
		X"A4",X"8D",X"3C",X"8D",X"24",X"34",X"02",X"D7",X"38",X"8E",X"C4",X"91",X"BD",X"FF",X"A4",X"96",
		X"39",X"8D",X"2C",X"8D",X"14",X"4D",X"27",X"04",X"0F",X"38",X"0F",X"39",X"AB",X"E0",X"19",X"C6",
		X"04",X"BD",X"CB",X"E6",X"BD",X"CC",X"0D",X"35",X"96",X"34",X"04",X"5D",X"26",X"03",X"4F",X"35",
		X"84",X"1E",X"89",X"86",X"99",X"8B",X"01",X"19",X"E0",X"E4",X"24",X"F9",X"EB",X"E0",X"39",X"34",
		X"02",X"1E",X"89",X"5F",X"4D",X"26",X"02",X"35",X"82",X"8B",X"99",X"19",X"5C",X"20",X"F5",X"34",
		X"36",X"8E",X"CE",X"CF",X"10",X"8E",X"C4",X"1D",X"C6",X"30",X"BD",X"CB",X"AF",X"8D",X"02",X"35",
		X"B6",X"34",X"36",X"10",X"8E",X"CE",X"CF",X"8E",X"B2",X"60",X"C6",X"30",X"A6",X"A0",X"BD",X"FF",
		X"AA",X"5A",X"26",X"F8",X"35",X"B6",X"CD",X"46",X"00",X"01",X"CD",X"51",X"00",X"05",X"CD",X"5E",
		X"00",X"09",X"CD",X"6A",X"00",X"0D",X"CD",X"75",X"00",X"11",X"CD",X"7F",X"00",X"15",X"CD",X"8A",
		X"00",X"19",X"CD",X"96",X"00",X"81",X"CD",X"A7",X"00",X"85",X"CD",X"B7",X"00",X"87",X"CD",X"C6",
		X"00",X"89",X"CD",X"D5",X"00",X"8B",X"CD",X"E6",X"00",X"8D",X"CD",X"F6",X"00",X"8F",X"CE",X"07",
		X"00",X"91",X"CE",X"17",X"00",X"93",X"CE",X"25",X"00",X"95",X"CE",X"2F",X"00",X"97",X"CE",X"3D",
		X"00",X"99",X"CE",X"4B",X"00",X"9B",X"CE",X"59",X"00",X"9D",X"CE",X"67",X"00",X"9F",X"CE",X"75",
		X"00",X"A1",X"CE",X"83",X"00",X"A3",X"CE",X"91",X"00",X"A5",X"CE",X"9F",X"00",X"A7",X"CE",X"AD",
		X"00",X"A9",X"CE",X"BC",X"00",X"7D",X"43",X"4F",X"49",X"4E",X"53",X"20",X"4C",X"45",X"46",X"54",
		X"2F",X"43",X"4F",X"49",X"4E",X"53",X"20",X"43",X"45",X"4E",X"54",X"45",X"52",X"2F",X"43",X"4F",
		X"49",X"4E",X"53",X"20",X"52",X"49",X"47",X"48",X"54",X"2F",X"54",X"4F",X"54",X"41",X"4C",X"20",
		X"50",X"41",X"49",X"44",X"2F",X"53",X"48",X"49",X"50",X"53",X"20",X"57",X"4F",X"4E",X"2F",X"54",
		X"4F",X"54",X"41",X"4C",X"20",X"54",X"49",X"4D",X"45",X"2F",X"54",X"4F",X"54",X"41",X"4C",X"20",
		X"53",X"48",X"49",X"50",X"53",X"2F",X"42",X"4F",X"4E",X"55",X"53",X"20",X"53",X"48",X"49",X"50",
		X"20",X"4C",X"45",X"56",X"45",X"4C",X"2F",X"4E",X"55",X"4D",X"42",X"45",X"52",X"20",X"4F",X"46",
		X"20",X"53",X"48",X"49",X"50",X"53",X"2F",X"43",X"4F",X"49",X"4E",X"41",X"47",X"45",X"20",X"53",
		X"45",X"4C",X"45",X"43",X"54",X"2F",X"4C",X"45",X"46",X"54",X"20",X"43",X"4F",X"49",X"4E",X"20",
		X"4D",X"55",X"4C",X"54",X"2F",X"43",X"45",X"4E",X"54",X"45",X"52",X"20",X"43",X"4F",X"49",X"4E",
		X"20",X"4D",X"55",X"4C",X"54",X"2F",X"52",X"49",X"47",X"48",X"54",X"20",X"43",X"4F",X"49",X"4E",
		X"20",X"4D",X"55",X"4C",X"54",X"2F",X"43",X"4F",X"49",X"4E",X"53",X"20",X"46",X"4F",X"52",X"20",
		X"43",X"52",X"45",X"44",X"49",X"54",X"2F",X"43",X"4F",X"49",X"4E",X"53",X"20",X"46",X"4F",X"52",
		X"20",X"42",X"4F",X"4E",X"55",X"53",X"2F",X"4D",X"49",X"4E",X"49",X"4D",X"55",X"4D",X"20",X"43",
		X"4F",X"49",X"4E",X"53",X"2F",X"46",X"52",X"45",X"45",X"20",X"50",X"4C",X"41",X"59",X"2F",X"47",
		X"41",X"4D",X"45",X"20",X"41",X"44",X"4A",X"55",X"53",X"54",X"20",X"31",X"2F",X"47",X"41",X"4D",
		X"45",X"20",X"41",X"44",X"4A",X"55",X"53",X"54",X"20",X"32",X"2F",X"47",X"41",X"4D",X"45",X"20",
		X"41",X"44",X"4A",X"55",X"53",X"54",X"20",X"33",X"2F",X"47",X"41",X"4D",X"45",X"20",X"41",X"44",
		X"4A",X"55",X"53",X"54",X"20",X"34",X"2F",X"47",X"41",X"4D",X"45",X"20",X"41",X"44",X"4A",X"55",
		X"53",X"54",X"20",X"35",X"2F",X"47",X"41",X"4D",X"45",X"20",X"41",X"44",X"4A",X"55",X"53",X"54",
		X"20",X"36",X"2F",X"47",X"41",X"4D",X"45",X"20",X"41",X"44",X"4A",X"55",X"53",X"54",X"20",X"37",
		X"2F",X"47",X"41",X"4D",X"45",X"20",X"41",X"44",X"4A",X"55",X"53",X"54",X"20",X"38",X"2F",X"47",
		X"41",X"4D",X"45",X"20",X"41",X"44",X"4A",X"55",X"53",X"54",X"20",X"39",X"2F",X"47",X"41",X"4D",
		X"45",X"20",X"41",X"44",X"4A",X"55",X"53",X"54",X"20",X"31",X"30",X"2F",X"53",X"50",X"45",X"43",
		X"49",X"41",X"4C",X"20",X"46",X"55",X"4E",X"43",X"54",X"49",X"4F",X"4E",X"2F",X"FF",X"FF",X"02",
		X"12",X"70",X"44",X"52",X"4A",X"01",X"83",X"15",X"53",X"41",X"4D",X"01",X"59",X"20",X"4C",X"45",
		X"44",X"01",X"42",X"85",X"50",X"47",X"44",X"01",X"25",X"20",X"43",X"52",X"42",X"01",X"10",X"35",
		X"4D",X"52",X"53",X"00",X"82",X"65",X"53",X"53",X"52",X"00",X"60",X"10",X"54",X"4D",X"48",X"00",
		X"5A",X"01",X"00",X"03",X"03",X"01",X"04",X"01",X"01",X"00",X"00",X"00",X"05",X"15",X"01",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"04",X"01",X"02",X"04",X"00",X"06",X"00",X"01",X"01",
		X"00",X"00",X"01",X"04",X"01",X"01",X"00",X"00",X"01",X"16",X"06",X"02",X"00",X"00",X"01",X"04",
		X"01",X"02",X"00",X"00",X"01",X"00",X"04",X"01",X"00",X"00",X"01",X"00",X"02",X"01",X"00",X"00",
		X"01",X"00",X"02",X"02",X"00",X"00",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",
		X"31",X"39",X"38",X"30",X"20",X"2D",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",
		X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"4A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"C0",X"15",X"7E",X"C0",X"92",X"7E",X"C2",X"62",X"7E",X"C2",X"9A",X"C4",X"50",X"7E",X"C5",
		X"D0",X"C6",X"BA",X"C7",X"72",X"DC",X"20",X"C4",X"E0",X"DD",X"17",X"C3",X"26",X"10",X"DD",X"15",
		X"0F",X"0F",X"8E",X"C3",X"4F",X"9F",X"09",X"86",X"E0",X"97",X"11",X"BD",X"C2",X"AA",X"8E",X"00",
		X"10",X"9C",X"15",X"27",X"12",X"96",X"0D",X"2A",X"04",X"0A",X"11",X"20",X"02",X"0C",X"11",X"BD",
		X"C2",X"AA",X"30",X"88",X"20",X"20",X"EA",X"DC",X"09",X"DD",X"03",X"96",X"0F",X"97",X"00",X"96",
		X"0D",X"97",X"01",X"96",X"11",X"97",X"02",X"8E",X"B7",X"00",X"9F",X"05",X"8E",X"BA",X"90",X"9F",
		X"07",X"DC",X"15",X"83",X"00",X"20",X"DD",X"15",X"10",X"93",X"17",X"2B",X"05",X"BD",X"C1",X"2C",
		X"20",X"EF",X"DC",X"03",X"DD",X"0B",X"96",X"00",X"97",X"10",X"96",X"01",X"97",X"0E",X"96",X"02",
		X"97",X"12",X"10",X"8E",X"BE",X"20",X"8E",X"00",X"00",X"AF",X"A1",X"10",X"8C",X"BF",X"50",X"26",
		X"F8",X"39",X"DC",X"20",X"C4",X"E0",X"93",X"15",X"58",X"49",X"58",X"49",X"58",X"49",X"97",X"00",
		X"27",X"20",X"2B",X"10",X"DC",X"15",X"C3",X"00",X"20",X"DD",X"15",X"BD",X"C1",X"CD",X"0A",X"00",
		X"26",X"F2",X"20",X"0E",X"DC",X"15",X"83",X"00",X"20",X"DD",X"15",X"BD",X"C1",X"2C",X"0C",X"00",
		X"26",X"F2",X"DC",X"20",X"C4",X"E0",X"DD",X"15",X"8E",X"00",X"00",X"10",X"8E",X"BE",X"20",X"10",
		X"DF",X"13",X"10",X"DE",X"05",X"C5",X"20",X"26",X"03",X"10",X"DE",X"07",X"86",X"98",X"AF",X"B4",
		X"35",X"44",X"ED",X"A4",X"EF",X"B1",X"4A",X"AF",X"B4",X"35",X"44",X"ED",X"A4",X"EF",X"B1",X"4A",
		X"AF",X"B4",X"35",X"44",X"ED",X"A4",X"EF",X"B1",X"4A",X"AF",X"B4",X"35",X"44",X"ED",X"A4",X"EF",
		X"B1",X"4A",X"AF",X"B4",X"35",X"44",X"ED",X"A4",X"EF",X"B1",X"4A",X"AF",X"B4",X"35",X"44",X"ED",
		X"A4",X"EF",X"B1",X"4A",X"AF",X"B4",X"35",X"44",X"ED",X"A4",X"EF",X"B1",X"4A",X"AF",X"B4",X"35",
		X"44",X"ED",X"A4",X"EF",X"B1",X"4A",X"26",X"B6",X"10",X"DE",X"13",X"39",X"BD",X"C3",X"23",X"2B",
		X"04",X"0A",X"12",X"20",X"02",X"0C",X"12",X"86",X"20",X"95",X"16",X"26",X"48",X"9E",X"07",X"BD",
		X"C2",X"F6",X"2B",X"20",X"0A",X"11",X"96",X"11",X"A7",X"84",X"A7",X"89",X"01",X"C8",X"CC",X"70",
		X"07",X"ED",X"01",X"ED",X"89",X"01",X"C9",X"30",X"03",X"8C",X"BC",X"58",X"26",X"03",X"8E",X"BA",
		X"90",X"9F",X"07",X"39",X"96",X"11",X"A7",X"84",X"A7",X"89",X"01",X"C8",X"4C",X"97",X"11",X"CC",
		X"07",X"70",X"ED",X"01",X"ED",X"89",X"01",X"C9",X"30",X"03",X"8C",X"BC",X"58",X"26",X"03",X"8E",
		X"BA",X"90",X"9F",X"07",X"39",X"9E",X"05",X"BD",X"C2",X"F6",X"2B",X"20",X"0A",X"11",X"96",X"11",
		X"A7",X"84",X"A7",X"89",X"01",X"C8",X"CC",X"70",X"07",X"ED",X"01",X"ED",X"89",X"01",X"C9",X"30",
		X"03",X"8C",X"B8",X"C8",X"26",X"03",X"8E",X"B7",X"00",X"9F",X"05",X"39",X"96",X"11",X"A7",X"84",
		X"A7",X"89",X"01",X"C8",X"4C",X"97",X"11",X"CC",X"07",X"70",X"ED",X"01",X"ED",X"89",X"01",X"C9",
		X"30",X"03",X"8C",X"B8",X"C8",X"26",X"03",X"8E",X"B7",X"00",X"9F",X"05",X"39",X"96",X"0D",X"2A",
		X"04",X"0A",X"11",X"20",X"02",X"0C",X"11",X"BD",X"C2",X"AA",X"86",X"20",X"95",X"16",X"27",X"41",
		X"9E",X"07",X"30",X"1D",X"8C",X"BA",X"8D",X"26",X"03",X"8E",X"BC",X"55",X"9F",X"07",X"96",X"0E",
		X"2A",X"17",X"0A",X"12",X"96",X"12",X"A7",X"84",X"A7",X"89",X"01",X"C8",X"CC",X"07",X"70",X"ED",
		X"01",X"ED",X"89",X"01",X"C9",X"BD",X"C2",X"D0",X"39",X"96",X"12",X"A7",X"84",X"A7",X"89",X"01",
		X"C8",X"4C",X"97",X"12",X"CC",X"70",X"07",X"ED",X"01",X"ED",X"89",X"01",X"C9",X"BD",X"C2",X"D0",
		X"39",X"9E",X"05",X"30",X"1D",X"8C",X"B6",X"FD",X"26",X"03",X"8E",X"B8",X"C5",X"9F",X"05",X"96",
		X"0E",X"2A",X"17",X"0A",X"12",X"96",X"12",X"A7",X"84",X"A7",X"89",X"01",X"C8",X"CC",X"07",X"70",
		X"ED",X"01",X"ED",X"89",X"01",X"C9",X"BD",X"C2",X"D0",X"39",X"96",X"12",X"A7",X"84",X"A7",X"89",
		X"01",X"C8",X"4C",X"97",X"12",X"CC",X"70",X"07",X"ED",X"01",X"ED",X"89",X"01",X"C9",X"BD",X"C2",
		X"D0",X"39",X"8E",X"C3",X"50",X"9F",X"0B",X"A6",X"84",X"97",X"0E",X"86",X"07",X"97",X"10",X"86",
		X"E0",X"97",X"12",X"8E",X"B3",X"00",X"96",X"12",X"A7",X"80",X"96",X"0E",X"2A",X"04",X"0A",X"12",
		X"20",X"02",X"0C",X"12",X"BD",X"C2",X"D0",X"96",X"0E",X"2A",X"04",X"0A",X"12",X"20",X"02",X"0C",
		X"12",X"BD",X"C2",X"D0",X"8C",X"B7",X"00",X"26",X"DD",X"39",X"8E",X"00",X"00",X"10",X"8E",X"BE",
		X"20",X"AF",X"B1",X"10",X"8C",X"BF",X"50",X"26",X"F8",X"39",X"96",X"0F",X"27",X"0A",X"0A",X"0F",
		X"96",X"0D",X"48",X"89",X"00",X"97",X"0D",X"39",X"DE",X"09",X"33",X"41",X"11",X"83",X"C4",X"50",
		X"26",X"03",X"CE",X"C3",X"50",X"DF",X"09",X"86",X"07",X"97",X"0F",X"A6",X"C4",X"97",X"0D",X"39",
		X"96",X"10",X"27",X"0A",X"0A",X"10",X"96",X"0E",X"48",X"89",X"00",X"97",X"0E",X"39",X"DE",X"0B",
		X"33",X"41",X"11",X"83",X"C4",X"50",X"26",X"03",X"CE",X"C3",X"50",X"DF",X"0B",X"86",X"07",X"97",
		X"10",X"A6",X"C4",X"97",X"0E",X"39",X"96",X"0F",X"81",X"07",X"27",X"0C",X"0C",X"0F",X"96",X"0D",
		X"44",X"24",X"02",X"8B",X"80",X"97",X"0D",X"39",X"DE",X"09",X"11",X"83",X"C3",X"50",X"26",X"03",
		X"CE",X"C4",X"50",X"33",X"5F",X"DF",X"09",X"0F",X"0F",X"A6",X"C4",X"44",X"24",X"02",X"8B",X"80",
		X"97",X"0D",X"39",X"96",X"10",X"81",X"07",X"27",X"0C",X"0C",X"10",X"96",X"0E",X"44",X"24",X"02",
		X"8B",X"80",X"97",X"0E",X"39",X"DE",X"0B",X"11",X"83",X"C3",X"50",X"26",X"03",X"CE",X"C4",X"50",
		X"33",X"5F",X"DF",X"0B",X"0F",X"10",X"A6",X"C4",X"44",X"24",X"02",X"8B",X"80",X"97",X"0E",X"39",
		X"2A",X"AA",X"AA",X"AA",X"AA",X"AA",X"AB",X"A1",X"D5",X"55",X"55",X"55",X"55",X"55",X"AA",X"BF",
		X"FF",X"FF",X"FF",X"C0",X"00",X"00",X"00",X"55",X"55",X"57",X"FF",X"C0",X"01",X"55",X"55",X"55",
		X"55",X"55",X"55",X"5F",X"E0",X"15",X"55",X"55",X"57",X"FF",X"F0",X"00",X"15",X"55",X"5F",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"05",X"55",X"7F",X"FF",X"E0",X"00",X"05",X"55",X"55",
		X"55",X"55",X"FC",X"05",X"55",X"55",X"50",X"01",X"FF",X"FF",X"FF",X"C0",X"00",X"0A",X"AA",X"AA",
		X"AA",X"FF",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"00",X"00",X"1F",X"E0",X"00",X"55",X"55",
		X"55",X"40",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"B5",X"57",X"AA",X"AA",X"AA",X"F5",X"7F",X"D5",
		X"55",X"55",X"57",X"FF",X"80",X"07",X"E0",X"7F",X"F1",X"55",X"7F",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"EF",X"76",X"91",X"11",X"11",X"5E",X"DB",X"E9",X"84",X"77",X"EC",X"C4",X"87",
		X"47",X"98",X"08",X"98",X"3F",X"C3",X"CB",X"DB",X"9F",X"C7",X"5F",X"2F",X"C7",X"7D",X"EF",X"BF",
		X"FA",X"4C",X"57",X"2B",X"61",X"EF",X"EF",X"FB",X"F7",X"E8",X"00",X"20",X"40",X"00",X"14",X"04",
		X"04",X"3C",X"06",X"00",X"1D",X"07",X"3C",X"E1",X"A5",X"55",X"55",X"45",X"2A",X"AA",X"AA",X"AA",
		X"A8",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"AA",X"AA",X"FE",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EA",X"AA",X"AA",X"A8",X"02",X"AA",X"AA",X"AA",X"AA",
		X"BF",X"BE",X"3E",X"63",X"FF",X"E0",X"D8",X"1C",X"18",X"2A",X"AB",X"1E",X"77",X"7A",X"AF",X"A8",
		X"40",X"70",X"7D",X"40",X"0B",X"FB",X"FA",X"FF",X"C1",X"53",X"54",X"75",X"70",X"03",X"00",X"00",
		X"25",X"70",X"07",X"26",X"77",X"00",X"26",X"07",X"70",X"24",X"07",X"70",X"23",X"07",X"70",X"23",
		X"70",X"07",X"24",X"07",X"70",X"25",X"70",X"07",X"26",X"77",X"00",X"25",X"07",X"70",X"24",X"07",
		X"70",X"23",X"07",X"70",X"21",X"07",X"70",X"22",X"70",X"07",X"24",X"77",X"00",X"24",X"70",X"07",
		X"26",X"77",X"00",X"26",X"77",X"00",X"25",X"77",X"00",X"25",X"70",X"07",X"26",X"77",X"00",X"24",
		X"07",X"70",X"23",X"70",X"07",X"25",X"77",X"00",X"26",X"70",X"07",X"26",X"77",X"00",X"26",X"77",
		X"00",X"25",X"07",X"70",X"23",X"07",X"70",X"22",X"07",X"70",X"21",X"77",X"00",X"21",X"70",X"07",
		X"23",X"70",X"07",X"25",X"70",X"07",X"25",X"07",X"70",X"25",X"77",X"00",X"25",X"77",X"00",X"24",
		X"77",X"00",X"22",X"07",X"70",X"20",X"07",X"70",X"1E",X"07",X"70",X"1C",X"07",X"70",X"1D",X"70",
		X"07",X"1F",X"70",X"07",X"21",X"70",X"07",X"22",X"70",X"07",X"24",X"70",X"07",X"26",X"70",X"07",
		X"26",X"77",X"00",X"26",X"77",X"00",X"26",X"77",X"00",X"26",X"77",X"00",X"26",X"77",X"00",X"25",
		X"77",X"00",X"25",X"70",X"07",X"26",X"77",X"00",X"24",X"07",X"70",X"23",X"77",X"00",X"24",X"77",
		X"00",X"22",X"07",X"70",X"23",X"70",X"07",X"22",X"07",X"70",X"21",X"70",X"07",X"23",X"70",X"07",
		X"25",X"70",X"07",X"26",X"77",X"00",X"26",X"07",X"70",X"24",X"07",X"70",X"23",X"07",X"70",X"23",
		X"70",X"07",X"24",X"07",X"70",X"25",X"70",X"07",X"26",X"77",X"00",X"25",X"07",X"70",X"24",X"07",
		X"70",X"23",X"07",X"70",X"21",X"07",X"70",X"22",X"70",X"07",X"24",X"77",X"00",X"24",X"70",X"07",
		X"26",X"77",X"00",X"26",X"77",X"00",X"25",X"77",X"00",X"25",X"70",X"07",X"26",X"77",X"00",X"24",
		X"07",X"70",X"23",X"70",X"07",X"25",X"77",X"00",X"26",X"70",X"07",X"26",X"77",X"00",X"26",X"77",
		X"00",X"25",X"07",X"70",X"23",X"07",X"70",X"22",X"07",X"70",X"21",X"77",X"00",X"21",X"70",X"07",
		X"23",X"70",X"07",X"25",X"70",X"07",X"25",X"07",X"70",X"25",X"77",X"00",X"25",X"77",X"00",X"24",
		X"77",X"00",X"22",X"07",X"70",X"20",X"07",X"70",X"1E",X"07",X"70",X"1C",X"07",X"70",X"1D",X"70",
		X"07",X"1F",X"70",X"07",X"21",X"70",X"07",X"22",X"70",X"07",X"24",X"70",X"07",X"26",X"70",X"07",
		X"26",X"77",X"00",X"26",X"77",X"00",X"26",X"77",X"00",X"26",X"77",X"00",X"26",X"77",X"00",X"25",
		X"77",X"00",X"25",X"70",X"07",X"26",X"77",X"00",X"24",X"07",X"70",X"23",X"77",X"00",X"24",X"77",
		X"00",X"22",X"07",X"70",X"23",X"70",X"07",X"22",X"07",X"70",X"21",X"70",X"07",X"23",X"70",X"07",
		X"35",X"06",X"ED",X"49",X"9F",X"00",X"CC",X"08",X"08",X"DD",X"04",X"CC",X"17",X"32",X"DD",X"06",
		X"10",X"8E",X"B3",X"00",X"96",X"00",X"5F",X"ED",X"22",X"96",X"01",X"ED",X"24",X"96",X"05",X"44",
		X"98",X"05",X"44",X"44",X"06",X"04",X"06",X"05",X"96",X"04",X"84",X"01",X"80",X"01",X"D6",X"05",
		X"ED",X"26",X"2A",X"02",X"43",X"53",X"34",X"06",X"96",X"07",X"44",X"98",X"07",X"44",X"44",X"06",
		X"06",X"06",X"07",X"96",X"06",X"84",X"03",X"80",X"02",X"D6",X"07",X"ED",X"28",X"2A",X"02",X"43",
		X"53",X"44",X"56",X"E3",X"E1",X"10",X"83",X"01",X"6A",X"24",X"B9",X"8E",X"00",X"00",X"AF",X"A4",
		X"31",X"2A",X"10",X"8C",X"B8",X"00",X"26",X"AC",X"8E",X"C6",X"AB",X"9F",X"02",X"86",X"38",X"97",
		X"01",X"86",X"01",X"8E",X"C6",X"49",X"7E",X"FF",X"D1",X"8E",X"00",X"00",X"10",X"8E",X"B3",X"00",
		X"A6",X"9F",X"A0",X"02",X"97",X"31",X"27",X"50",X"EE",X"A4",X"AF",X"C4",X"AF",X"C9",X"01",X"00",
		X"EC",X"28",X"E3",X"24",X"81",X"2A",X"25",X"28",X"ED",X"24",X"A7",X"21",X"EC",X"26",X"E3",X"22",
		X"81",X"98",X"22",X"1C",X"ED",X"22",X"A7",X"A4",X"5D",X"2B",X"07",X"CC",X"BB",X"BB",X"ED",X"B4",
		X"20",X"0E",X"EE",X"A4",X"CC",X"0B",X"0B",X"ED",X"C4",X"CC",X"B0",X"B0",X"ED",X"C9",X"01",X"00",
		X"31",X"2A",X"10",X"8C",X"B8",X"00",X"26",X"C0",X"0A",X"01",X"26",X"A5",X"DE",X"02",X"33",X"41",
		X"DF",X"02",X"86",X"04",X"97",X"01",X"20",X"99",X"6E",X"D8",X"09",X"FF",X"7F",X"3F",X"37",X"2F",
		X"27",X"1F",X"17",X"07",X"06",X"05",X"04",X"03",X"02",X"00",X"14",X"00",X"00",X"00",X"0F",X"14",
		X"14",X"14",X"03",X"00",X"00",X"00",X"00",X"03",X"04",X"05",X"06",X"00",X"00",X"00",X"00",X"01",
		X"03",X"04",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"1E",X"00",X"00",X"00",X"1E",X"19",X"14",X"10",X"05",X"00",X"00",X"00",X"05",X"05",
		X"05",X"05",X"60",X"00",X"03",X"02",X"16",X"1E",X"26",X"2E",X"01",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"FF",X"00",X"10",X"00",X"70",X"B0",X"00",X"00",X"80",X"10",X"FC",X"FE",X"4A",X"3A",
		X"2A",X"2A",X"30",X"00",X"00",X"00",X"20",X"28",X"2C",X"30",X"02",X"00",X"00",X"00",X"01",X"01",
		X"02",X"02",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"FF",X"00",X"08",X"06",X"62",X"E0",
		X"02",X"12",X"60",X"00",X"08",X"04",X"0C",X"1C",X"24",X"28",X"FF",X"08",X"FE",X"FE",X"2A",X"22",
		X"1E",X"1C",X"60",X"00",X"08",X"02",X"16",X"1E",X"20",X"22",X"28",X"0A",X"FE",X"FF",X"19",X"19",
		X"19",X"19",X"3F",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"3F",X"C0",X"18",X"F4",X"FC",X"D4",X"C4",
		X"A4",X"94",X"0A",X"03",X"FF",X"FF",X"0F",X"0D",X"0C",X"0A",X"C8",X"28",X"F4",X"F8",X"F0",X"DC",
		X"C8",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"8E",X"C0",X"0C",X"7E",X"C0",X"36",X"C6",
		X"28",X"20",X"F1",X"C6",X"80",X"20",X"ED",X"10",X"8E",X"C9",X"FE",X"BD",X"CA",X"97",X"7E",X"CB",
		X"3B",X"C6",X"A5",X"8E",X"C0",X"01",X"7E",X"C0",X"36",X"BD",X"CA",X"69",X"BD",X"CA",X"2A",X"8D",
		X"F0",X"CE",X"C0",X"D7",X"8E",X"28",X"20",X"BD",X"CA",X"69",X"BD",X"C0",X"3C",X"10",X"8E",X"C0",
		X"61",X"BD",X"C0",X"6D",X"10",X"8E",X"05",X"DC",X"BD",X"CA",X"44",X"0D",X"49",X"26",X"60",X"0F",
		X"3C",X"86",X"01",X"97",X"3B",X"32",X"E8",X"E0",X"BD",X"FF",X"BC",X"CE",X"C0",X"D7",X"8E",X"28",
		X"20",X"BD",X"CA",X"69",X"BD",X"C0",X"3C",X"0F",X"3A",X"10",X"8E",X"C0",X"65",X"BD",X"C0",X"66",
		X"BD",X"CA",X"69",X"86",X"20",X"1F",X"89",X"5A",X"30",X"E4",X"A7",X"80",X"5A",X"26",X"FB",X"86",
		X"17",X"A7",X"80",X"30",X"E4",X"BD",X"CA",X"57",X"8E",X"CC",X"00",X"BD",X"C0",X"39",X"C5",X"02");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
